// soc_system.v

// Generated using ACDS version 22.1 917

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        aes_reset_in_reset,      //      aes_reset_in.reset
		output wire [31:0] aes_reset_out_export,    //     aes_reset_out.export
		input  wire        clk_clk,                 //               clk.clk
		input  wire [31:0] locked_phi_in_export,    //     locked_phi_in.export
		output wire        locked_phi_out_export,   //    locked_phi_out.export
		input  wire [31:0] locked_theta_in_export,  //   locked_theta_in.export
		output wire        locked_theta_out_export, //  locked_theta_out.export
		output wire [14:0] memory_mem_a,            //            memory.mem_a
		output wire [2:0]  memory_mem_ba,           //                  .mem_ba
		output wire        memory_mem_ck,           //                  .mem_ck
		output wire        memory_mem_ck_n,         //                  .mem_ck_n
		output wire        memory_mem_cke,          //                  .mem_cke
		output wire        memory_mem_cs_n,         //                  .mem_cs_n
		output wire        memory_mem_ras_n,        //                  .mem_ras_n
		output wire        memory_mem_cas_n,        //                  .mem_cas_n
		output wire        memory_mem_we_n,         //                  .mem_we_n
		output wire        memory_mem_reset_n,      //                  .mem_reset_n
		inout  wire [31:0] memory_mem_dq,           //                  .mem_dq
		inout  wire [3:0]  memory_mem_dqs,          //                  .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,        //                  .mem_dqs_n
		output wire        memory_mem_odt,          //                  .mem_odt
		output wire [3:0]  memory_mem_dm,           //                  .mem_dm
		input  wire        memory_oct_rzqin,        //                  .oct_rzqin
		input  wire        reset_phi_in_reset,      //      reset_phi_in.reset
		output wire [31:0] reset_phi_out_export,    //     reset_phi_out.export
		input  wire        reset_theta_in_reset,    //    reset_theta_in.reset
		output wire [31:0] reset_theta_out_export,  //   reset_theta_out.export
		input  wire        tdc_reset_in_reset,      //      tdc_reset_in.reset
		output wire [31:0] tdc_reset_out_export,    //     tdc_reset_out.export
		input  wire        theta_clks_refclk_clk    // theta_clks_refclk.clk
	);

	wire          pulsegenerator_avalon_streaming_source_valid;                       // pulsegenerator:M_AVST_VALID -> tdc_0:S_AVST_VALID
	wire    [7:0] pulsegenerator_avalon_streaming_source_data;                        // pulsegenerator:M_AVST_DATA -> tdc_0:S_AVST_DATA
	wire          pulsegenerator_avalon_streaming_source_ready;                       // tdc_0:S_AVST_READY -> pulsegenerator:M_AVST_READY
	wire          tdc_0_avalon_streaming_source_valid;                                // tdc_0:M_AVST_VALID -> tdc_to_dma_dc_fifo:in_valid
	wire  [255:0] tdc_0_avalon_streaming_source_data;                                 // tdc_0:M_AVST_DATA -> tdc_to_dma_dc_fifo:in_data
	wire          tdc_0_avalon_streaming_source_ready;                                // tdc_to_dma_dc_fifo:in_ready -> tdc_0:M_AVST_READY
	wire          ip_sync_avalon_streaming_source_valid;                              // ip_sync:M_AVST_VALID -> ip_sync_to_pulsegenerator_cdc:in_valid
	wire    [7:0] ip_sync_avalon_streaming_source_data;                               // ip_sync:M_AVST_DATA -> ip_sync_to_pulsegenerator_cdc:in_data
	wire          ip_sync_avalon_streaming_source_ready;                              // ip_sync_to_pulsegenerator_cdc:in_ready -> ip_sync:M_AVST_READY
	wire          ip_sync_to_pulsegenerator_cdc_out_valid;                            // ip_sync_to_pulsegenerator_cdc:out_valid -> pulsegenerator:S_AVST_VALID
	wire    [7:0] ip_sync_to_pulsegenerator_cdc_out_data;                             // ip_sync_to_pulsegenerator_cdc:out_data -> pulsegenerator:S_AVST_DATA
	wire          ip_sync_to_pulsegenerator_cdc_out_ready;                            // pulsegenerator:S_AVST_READY -> ip_sync_to_pulsegenerator_cdc:out_ready
	wire          tdc_to_dma_dc_fifo_out_valid;                                       // tdc_to_dma_dc_fifo:out_valid -> DMA_to_SDRAM:st_sink_valid
	wire  [255:0] tdc_to_dma_dc_fifo_out_data;                                        // tdc_to_dma_dc_fifo:out_data -> DMA_to_SDRAM:st_sink_data
	wire          tdc_to_dma_dc_fifo_out_ready;                                       // DMA_to_SDRAM:st_sink_ready -> tdc_to_dma_dc_fifo:out_ready
	wire          theta_clks_outclk0_clk;                                             // theta_clks:outclk_0 -> [ip_sync_to_pulsegenerator_cdc:out_clk, mm_interconnect_3:theta_clks_outclk0_clk, pulsegenerator:S_AXI_ACLK, pulsegenerator_cdc:m0_clk, reset_bridge_launch:clk, rst_controller_003:clk, rst_controller_006:clk, tdc_0:clk_launch]
	wire          shell_pll_outclk0_clk;                                              // shell_pll:outclk_0 -> [DMA_to_SDRAM:clock_clk, aes_reset_pio:clk, hps_0:f2h_sdram0_clk, hps_0:h2f_axi_clk, hps_0:h2f_lw_axi_clk, ipsync_bridge:s0_clk, mm_interconnect_1:shell_pll_outclk0_clk, mm_interconnect_2:shell_pll_outclk0_clk, mm_interconnect_8:shell_pll_outclk0_clk, phi_locked:clk, phi_pll_reconfig_cdc:s0_clk, phi_pll_reset_pio:clk, pulsegenerator_cdc:s0_clk, reset_bridge_shell:clk, reset_bridge_tdc:clk, rst_controller:clk, rst_controller_007:clk, rst_controller_010:clk, tdc_reset_pio:clk, tdc_to_dma_dc_fifo:out_clk, theta_locked:clk, theta_pll_reconfig_cdc:s0_clk, theta_pll_reset_bridge:clk, theta_pll_reset_pio:clk]
	wire          theta_clks_outclk1_clk;                                             // theta_clks:outclk_1 -> [reset_bridge_capt:clk, rst_controller_008:clk, tdc_0:clk_capt, tdc_to_dma_dc_fifo:in_clk]
	wire          shell_pll_outclk1_clk;                                              // shell_pll:outclk_1 -> [aes:clk, aes_reset_controller:clk, ip_sync:clk, ip_sync_to_pulsegenerator_cdc:in_clk, ipsync_bridge:m0_clk, ipsync_to_aes_delay:m0_clk, ipsync_to_aes_delay:s0_clk, mm_interconnect_0:shell_pll_outclk1_clk, mm_interconnect_4:shell_pll_outclk1_clk, mm_interconnect_5:shell_pll_outclk1_clk, rst_controller_001:clk, rst_controller_002:clk]
	wire          phi_clk_cascade_out_export;                                         // phi_clk:cascade_out -> theta_clks:adjpllin
	wire   [63:0] theta_clks_reconfig_from_pll_reconfig_from_pll;                     // theta_clks:reconfig_from_pll -> theta_pll_reconfig:reconfig_from_pll
	wire   [63:0] phi_clk_reconfig_from_pll_reconfig_from_pll;                        // phi_clk:reconfig_from_pll -> phi_pll_reconfig:reconfig_from_pll
	wire   [63:0] theta_pll_reconfig_reconfig_to_pll_reconfig_to_pll;                 // theta_pll_reconfig:reconfig_to_pll -> theta_clks:reconfig_to_pll
	wire   [63:0] phi_pll_reconfig_reconfig_to_pll_reconfig_to_pll;                   // phi_pll_reconfig:reconfig_to_pll -> phi_clk:reconfig_to_pll
	wire          hps_0_h2f_reset_reset;                                              // hps_0:h2f_rst_n -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in0, rst_controller_002:reset_in1, rst_controller_003:reset_in0, rst_controller_003:reset_in1, rst_controller_004:reset_in0, rst_controller_004:reset_in1, rst_controller_005:reset_in0, rst_controller_005:reset_in1, rst_controller_006:reset_in0, rst_controller_006:reset_in1, rst_controller_007:reset_in0, rst_controller_007:reset_in1, rst_controller_008:reset_in0, rst_controller_008:reset_in1, rst_controller_009:reset_in0, rst_controller_009:reset_in1, rst_controller_010:reset_in0, shell_pll:rst]
	wire          reset_bridge_tdc_reset_out_reset;                                   // reset_bridge_tdc:reset_out -> [reset_bridge_capt:reset_in0, reset_bridge_launch:reset_in0, reset_bridge_shell:reset_in0]
	wire   [31:0] ip_sync_avalon_master_readdata;                                     // mm_interconnect_0:ip_sync_avalon_master_readdata -> ip_sync:M_AVMM_RDATA
	wire          ip_sync_avalon_master_waitrequest;                                  // mm_interconnect_0:ip_sync_avalon_master_waitrequest -> ip_sync:M_AVMM_WAITREQUEST
	wire    [7:0] ip_sync_avalon_master_address;                                      // ip_sync:M_AVMM_ADDR -> mm_interconnect_0:ip_sync_avalon_master_address
	wire    [3:0] ip_sync_avalon_master_byteenable;                                   // ip_sync:M_AVMM_BYTEENABLE -> mm_interconnect_0:ip_sync_avalon_master_byteenable
	wire          ip_sync_avalon_master_read;                                         // ip_sync:M_AVMM_R -> mm_interconnect_0:ip_sync_avalon_master_read
	wire          ip_sync_avalon_master_readdatavalid;                                // mm_interconnect_0:ip_sync_avalon_master_readdatavalid -> ip_sync:M_AVMM_READATAVALID
	wire          ip_sync_avalon_master_write;                                        // ip_sync:M_AVMM_W -> mm_interconnect_0:ip_sync_avalon_master_write
	wire   [31:0] ip_sync_avalon_master_writedata;                                    // ip_sync:M_AVMM_WDATA -> mm_interconnect_0:ip_sync_avalon_master_writedata
	wire          ip_sync_avalon_master_burstcount;                                   // ip_sync:M_AVMM_BURSTCOUNT -> mm_interconnect_0:ip_sync_avalon_master_burstcount
	wire   [31:0] mm_interconnect_0_ipsync_to_aes_delay_s0_readdata;                  // ipsync_to_aes_delay:s0_readdata -> mm_interconnect_0:ipsync_to_aes_delay_s0_readdata
	wire          mm_interconnect_0_ipsync_to_aes_delay_s0_waitrequest;               // ipsync_to_aes_delay:s0_waitrequest -> mm_interconnect_0:ipsync_to_aes_delay_s0_waitrequest
	wire          mm_interconnect_0_ipsync_to_aes_delay_s0_debugaccess;               // mm_interconnect_0:ipsync_to_aes_delay_s0_debugaccess -> ipsync_to_aes_delay:s0_debugaccess
	wire    [9:0] mm_interconnect_0_ipsync_to_aes_delay_s0_address;                   // mm_interconnect_0:ipsync_to_aes_delay_s0_address -> ipsync_to_aes_delay:s0_address
	wire          mm_interconnect_0_ipsync_to_aes_delay_s0_read;                      // mm_interconnect_0:ipsync_to_aes_delay_s0_read -> ipsync_to_aes_delay:s0_read
	wire    [3:0] mm_interconnect_0_ipsync_to_aes_delay_s0_byteenable;                // mm_interconnect_0:ipsync_to_aes_delay_s0_byteenable -> ipsync_to_aes_delay:s0_byteenable
	wire          mm_interconnect_0_ipsync_to_aes_delay_s0_readdatavalid;             // ipsync_to_aes_delay:s0_readdatavalid -> mm_interconnect_0:ipsync_to_aes_delay_s0_readdatavalid
	wire          mm_interconnect_0_ipsync_to_aes_delay_s0_write;                     // mm_interconnect_0:ipsync_to_aes_delay_s0_write -> ipsync_to_aes_delay:s0_write
	wire   [31:0] mm_interconnect_0_ipsync_to_aes_delay_s0_writedata;                 // mm_interconnect_0:ipsync_to_aes_delay_s0_writedata -> ipsync_to_aes_delay:s0_writedata
	wire    [0:0] mm_interconnect_0_ipsync_to_aes_delay_s0_burstcount;                // mm_interconnect_0:ipsync_to_aes_delay_s0_burstcount -> ipsync_to_aes_delay:s0_burstcount
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                       // hps_0:h2f_AWBURST -> mm_interconnect_1:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                         // hps_0:h2f_ARLEN -> mm_interconnect_1:hps_0_h2f_axi_master_arlen
	wire    [3:0] hps_0_h2f_axi_master_wstrb;                                         // hps_0:h2f_WSTRB -> mm_interconnect_1:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                        // mm_interconnect_1:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                           // mm_interconnect_1:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                        // hps_0:h2f_RREADY -> mm_interconnect_1:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                         // hps_0:h2f_AWLEN -> mm_interconnect_1:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                           // hps_0:h2f_WID -> mm_interconnect_1:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                       // hps_0:h2f_ARCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                        // hps_0:h2f_WVALID -> mm_interconnect_1:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                        // hps_0:h2f_ARADDR -> mm_interconnect_1:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                        // hps_0:h2f_ARPROT -> mm_interconnect_1:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                        // hps_0:h2f_AWPROT -> mm_interconnect_1:hps_0_h2f_axi_master_awprot
	wire   [31:0] hps_0_h2f_axi_master_wdata;                                         // hps_0:h2f_WDATA -> mm_interconnect_1:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                       // hps_0:h2f_ARVALID -> mm_interconnect_1:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                       // hps_0:h2f_AWCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                          // hps_0:h2f_ARID -> mm_interconnect_1:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                        // hps_0:h2f_ARLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                        // hps_0:h2f_AWLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                        // hps_0:h2f_AWADDR -> mm_interconnect_1:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                         // mm_interconnect_1:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                       // mm_interconnect_1:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire   [31:0] hps_0_h2f_axi_master_rdata;                                         // mm_interconnect_1:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                       // mm_interconnect_1:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                       // hps_0:h2f_ARBURST -> mm_interconnect_1:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                        // hps_0:h2f_ARSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                        // hps_0:h2f_BREADY -> mm_interconnect_1:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                         // mm_interconnect_1:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                         // hps_0:h2f_WLAST -> mm_interconnect_1:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                         // mm_interconnect_1:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                          // hps_0:h2f_AWID -> mm_interconnect_1:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                           // mm_interconnect_1:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                        // mm_interconnect_1:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                        // hps_0:h2f_AWSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                       // hps_0:h2f_AWVALID -> mm_interconnect_1:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                        // mm_interconnect_1:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire   [31:0] mm_interconnect_1_theta_pll_reconfig_cdc_s0_readdata;               // theta_pll_reconfig_cdc:s0_readdata -> mm_interconnect_1:theta_pll_reconfig_cdc_s0_readdata
	wire          mm_interconnect_1_theta_pll_reconfig_cdc_s0_waitrequest;            // theta_pll_reconfig_cdc:s0_waitrequest -> mm_interconnect_1:theta_pll_reconfig_cdc_s0_waitrequest
	wire          mm_interconnect_1_theta_pll_reconfig_cdc_s0_debugaccess;            // mm_interconnect_1:theta_pll_reconfig_cdc_s0_debugaccess -> theta_pll_reconfig_cdc:s0_debugaccess
	wire    [7:0] mm_interconnect_1_theta_pll_reconfig_cdc_s0_address;                // mm_interconnect_1:theta_pll_reconfig_cdc_s0_address -> theta_pll_reconfig_cdc:s0_address
	wire          mm_interconnect_1_theta_pll_reconfig_cdc_s0_read;                   // mm_interconnect_1:theta_pll_reconfig_cdc_s0_read -> theta_pll_reconfig_cdc:s0_read
	wire    [3:0] mm_interconnect_1_theta_pll_reconfig_cdc_s0_byteenable;             // mm_interconnect_1:theta_pll_reconfig_cdc_s0_byteenable -> theta_pll_reconfig_cdc:s0_byteenable
	wire          mm_interconnect_1_theta_pll_reconfig_cdc_s0_readdatavalid;          // theta_pll_reconfig_cdc:s0_readdatavalid -> mm_interconnect_1:theta_pll_reconfig_cdc_s0_readdatavalid
	wire          mm_interconnect_1_theta_pll_reconfig_cdc_s0_write;                  // mm_interconnect_1:theta_pll_reconfig_cdc_s0_write -> theta_pll_reconfig_cdc:s0_write
	wire   [31:0] mm_interconnect_1_theta_pll_reconfig_cdc_s0_writedata;              // mm_interconnect_1:theta_pll_reconfig_cdc_s0_writedata -> theta_pll_reconfig_cdc:s0_writedata
	wire    [0:0] mm_interconnect_1_theta_pll_reconfig_cdc_s0_burstcount;             // mm_interconnect_1:theta_pll_reconfig_cdc_s0_burstcount -> theta_pll_reconfig_cdc:s0_burstcount
	wire   [31:0] mm_interconnect_1_phi_pll_reconfig_cdc_s0_readdata;                 // phi_pll_reconfig_cdc:s0_readdata -> mm_interconnect_1:phi_pll_reconfig_cdc_s0_readdata
	wire          mm_interconnect_1_phi_pll_reconfig_cdc_s0_waitrequest;              // phi_pll_reconfig_cdc:s0_waitrequest -> mm_interconnect_1:phi_pll_reconfig_cdc_s0_waitrequest
	wire          mm_interconnect_1_phi_pll_reconfig_cdc_s0_debugaccess;              // mm_interconnect_1:phi_pll_reconfig_cdc_s0_debugaccess -> phi_pll_reconfig_cdc:s0_debugaccess
	wire    [7:0] mm_interconnect_1_phi_pll_reconfig_cdc_s0_address;                  // mm_interconnect_1:phi_pll_reconfig_cdc_s0_address -> phi_pll_reconfig_cdc:s0_address
	wire          mm_interconnect_1_phi_pll_reconfig_cdc_s0_read;                     // mm_interconnect_1:phi_pll_reconfig_cdc_s0_read -> phi_pll_reconfig_cdc:s0_read
	wire    [3:0] mm_interconnect_1_phi_pll_reconfig_cdc_s0_byteenable;               // mm_interconnect_1:phi_pll_reconfig_cdc_s0_byteenable -> phi_pll_reconfig_cdc:s0_byteenable
	wire          mm_interconnect_1_phi_pll_reconfig_cdc_s0_readdatavalid;            // phi_pll_reconfig_cdc:s0_readdatavalid -> mm_interconnect_1:phi_pll_reconfig_cdc_s0_readdatavalid
	wire          mm_interconnect_1_phi_pll_reconfig_cdc_s0_write;                    // mm_interconnect_1:phi_pll_reconfig_cdc_s0_write -> phi_pll_reconfig_cdc:s0_write
	wire   [31:0] mm_interconnect_1_phi_pll_reconfig_cdc_s0_writedata;                // mm_interconnect_1:phi_pll_reconfig_cdc_s0_writedata -> phi_pll_reconfig_cdc:s0_writedata
	wire    [0:0] mm_interconnect_1_phi_pll_reconfig_cdc_s0_burstcount;               // mm_interconnect_1:phi_pll_reconfig_cdc_s0_burstcount -> phi_pll_reconfig_cdc:s0_burstcount
	wire   [31:0] mm_interconnect_1_pulsegenerator_cdc_s0_readdata;                   // pulsegenerator_cdc:s0_readdata -> mm_interconnect_1:pulsegenerator_cdc_s0_readdata
	wire          mm_interconnect_1_pulsegenerator_cdc_s0_waitrequest;                // pulsegenerator_cdc:s0_waitrequest -> mm_interconnect_1:pulsegenerator_cdc_s0_waitrequest
	wire          mm_interconnect_1_pulsegenerator_cdc_s0_debugaccess;                // mm_interconnect_1:pulsegenerator_cdc_s0_debugaccess -> pulsegenerator_cdc:s0_debugaccess
	wire    [3:0] mm_interconnect_1_pulsegenerator_cdc_s0_address;                    // mm_interconnect_1:pulsegenerator_cdc_s0_address -> pulsegenerator_cdc:s0_address
	wire          mm_interconnect_1_pulsegenerator_cdc_s0_read;                       // mm_interconnect_1:pulsegenerator_cdc_s0_read -> pulsegenerator_cdc:s0_read
	wire    [3:0] mm_interconnect_1_pulsegenerator_cdc_s0_byteenable;                 // mm_interconnect_1:pulsegenerator_cdc_s0_byteenable -> pulsegenerator_cdc:s0_byteenable
	wire          mm_interconnect_1_pulsegenerator_cdc_s0_readdatavalid;              // pulsegenerator_cdc:s0_readdatavalid -> mm_interconnect_1:pulsegenerator_cdc_s0_readdatavalid
	wire          mm_interconnect_1_pulsegenerator_cdc_s0_write;                      // mm_interconnect_1:pulsegenerator_cdc_s0_write -> pulsegenerator_cdc:s0_write
	wire   [31:0] mm_interconnect_1_pulsegenerator_cdc_s0_writedata;                  // mm_interconnect_1:pulsegenerator_cdc_s0_writedata -> pulsegenerator_cdc:s0_writedata
	wire    [0:0] mm_interconnect_1_pulsegenerator_cdc_s0_burstcount;                 // mm_interconnect_1:pulsegenerator_cdc_s0_burstcount -> pulsegenerator_cdc:s0_burstcount
	wire   [31:0] mm_interconnect_1_ipsync_bridge_s0_readdata;                        // ipsync_bridge:s0_readdata -> mm_interconnect_1:ipsync_bridge_s0_readdata
	wire          mm_interconnect_1_ipsync_bridge_s0_waitrequest;                     // ipsync_bridge:s0_waitrequest -> mm_interconnect_1:ipsync_bridge_s0_waitrequest
	wire          mm_interconnect_1_ipsync_bridge_s0_debugaccess;                     // mm_interconnect_1:ipsync_bridge_s0_debugaccess -> ipsync_bridge:s0_debugaccess
	wire    [9:0] mm_interconnect_1_ipsync_bridge_s0_address;                         // mm_interconnect_1:ipsync_bridge_s0_address -> ipsync_bridge:s0_address
	wire          mm_interconnect_1_ipsync_bridge_s0_read;                            // mm_interconnect_1:ipsync_bridge_s0_read -> ipsync_bridge:s0_read
	wire    [3:0] mm_interconnect_1_ipsync_bridge_s0_byteenable;                      // mm_interconnect_1:ipsync_bridge_s0_byteenable -> ipsync_bridge:s0_byteenable
	wire          mm_interconnect_1_ipsync_bridge_s0_readdatavalid;                   // ipsync_bridge:s0_readdatavalid -> mm_interconnect_1:ipsync_bridge_s0_readdatavalid
	wire          mm_interconnect_1_ipsync_bridge_s0_write;                           // mm_interconnect_1:ipsync_bridge_s0_write -> ipsync_bridge:s0_write
	wire   [31:0] mm_interconnect_1_ipsync_bridge_s0_writedata;                       // mm_interconnect_1:ipsync_bridge_s0_writedata -> ipsync_bridge:s0_writedata
	wire    [0:0] mm_interconnect_1_ipsync_bridge_s0_burstcount;                      // mm_interconnect_1:ipsync_bridge_s0_burstcount -> ipsync_bridge:s0_burstcount
	wire          mm_interconnect_1_theta_pll_reset_pio_s1_chipselect;                // mm_interconnect_1:theta_pll_reset_pio_s1_chipselect -> theta_pll_reset_pio:chipselect
	wire   [31:0] mm_interconnect_1_theta_pll_reset_pio_s1_readdata;                  // theta_pll_reset_pio:readdata -> mm_interconnect_1:theta_pll_reset_pio_s1_readdata
	wire    [1:0] mm_interconnect_1_theta_pll_reset_pio_s1_address;                   // mm_interconnect_1:theta_pll_reset_pio_s1_address -> theta_pll_reset_pio:address
	wire          mm_interconnect_1_theta_pll_reset_pio_s1_write;                     // mm_interconnect_1:theta_pll_reset_pio_s1_write -> theta_pll_reset_pio:write_n
	wire   [31:0] mm_interconnect_1_theta_pll_reset_pio_s1_writedata;                 // mm_interconnect_1:theta_pll_reset_pio_s1_writedata -> theta_pll_reset_pio:writedata
	wire   [31:0] mm_interconnect_1_theta_locked_s1_readdata;                         // theta_locked:readdata -> mm_interconnect_1:theta_locked_s1_readdata
	wire    [1:0] mm_interconnect_1_theta_locked_s1_address;                          // mm_interconnect_1:theta_locked_s1_address -> theta_locked:address
	wire          mm_interconnect_1_phi_pll_reset_pio_s1_chipselect;                  // mm_interconnect_1:phi_pll_reset_pio_s1_chipselect -> phi_pll_reset_pio:chipselect
	wire   [31:0] mm_interconnect_1_phi_pll_reset_pio_s1_readdata;                    // phi_pll_reset_pio:readdata -> mm_interconnect_1:phi_pll_reset_pio_s1_readdata
	wire    [1:0] mm_interconnect_1_phi_pll_reset_pio_s1_address;                     // mm_interconnect_1:phi_pll_reset_pio_s1_address -> phi_pll_reset_pio:address
	wire          mm_interconnect_1_phi_pll_reset_pio_s1_write;                       // mm_interconnect_1:phi_pll_reset_pio_s1_write -> phi_pll_reset_pio:write_n
	wire   [31:0] mm_interconnect_1_phi_pll_reset_pio_s1_writedata;                   // mm_interconnect_1:phi_pll_reset_pio_s1_writedata -> phi_pll_reset_pio:writedata
	wire   [31:0] mm_interconnect_1_phi_locked_s1_readdata;                           // phi_locked:readdata -> mm_interconnect_1:phi_locked_s1_readdata
	wire    [1:0] mm_interconnect_1_phi_locked_s1_address;                            // mm_interconnect_1:phi_locked_s1_address -> phi_locked:address
	wire          mm_interconnect_1_tdc_reset_pio_s1_chipselect;                      // mm_interconnect_1:tdc_reset_pio_s1_chipselect -> tdc_reset_pio:chipselect
	wire   [31:0] mm_interconnect_1_tdc_reset_pio_s1_readdata;                        // tdc_reset_pio:readdata -> mm_interconnect_1:tdc_reset_pio_s1_readdata
	wire    [1:0] mm_interconnect_1_tdc_reset_pio_s1_address;                         // mm_interconnect_1:tdc_reset_pio_s1_address -> tdc_reset_pio:address
	wire          mm_interconnect_1_tdc_reset_pio_s1_write;                           // mm_interconnect_1:tdc_reset_pio_s1_write -> tdc_reset_pio:write_n
	wire   [31:0] mm_interconnect_1_tdc_reset_pio_s1_writedata;                       // mm_interconnect_1:tdc_reset_pio_s1_writedata -> tdc_reset_pio:writedata
	wire          mm_interconnect_1_aes_reset_pio_s1_chipselect;                      // mm_interconnect_1:aes_reset_pio_s1_chipselect -> aes_reset_pio:chipselect
	wire   [31:0] mm_interconnect_1_aes_reset_pio_s1_readdata;                        // aes_reset_pio:readdata -> mm_interconnect_1:aes_reset_pio_s1_readdata
	wire    [1:0] mm_interconnect_1_aes_reset_pio_s1_address;                         // mm_interconnect_1:aes_reset_pio_s1_address -> aes_reset_pio:address
	wire          mm_interconnect_1_aes_reset_pio_s1_write;                           // mm_interconnect_1:aes_reset_pio_s1_write -> aes_reset_pio:write_n
	wire   [31:0] mm_interconnect_1_aes_reset_pio_s1_writedata;                       // mm_interconnect_1:aes_reset_pio_s1_writedata -> aes_reset_pio:writedata
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                    // hps_0:h2f_lw_AWBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                      // hps_0:h2f_lw_ARLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                      // hps_0:h2f_lw_WSTRB -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                                     // mm_interconnect_2:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                        // mm_interconnect_2:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                                     // hps_0:h2f_lw_RREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                      // hps_0:h2f_lw_AWLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                        // hps_0:h2f_lw_WID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                    // hps_0:h2f_lw_ARCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                                     // hps_0:h2f_lw_WVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                     // hps_0:h2f_lw_ARADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                     // hps_0:h2f_lw_ARPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                     // hps_0:h2f_lw_AWPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                      // hps_0:h2f_lw_WDATA -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                                    // hps_0:h2f_lw_ARVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                    // hps_0:h2f_lw_AWCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                       // hps_0:h2f_lw_ARID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                     // hps_0:h2f_lw_ARLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                     // hps_0:h2f_lw_AWLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                     // hps_0:h2f_lw_AWADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                      // mm_interconnect_2:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                                    // mm_interconnect_2:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                      // mm_interconnect_2:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                                    // mm_interconnect_2:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                    // hps_0:h2f_lw_ARBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                     // hps_0:h2f_lw_ARSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                                     // hps_0:h2f_lw_BREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                                      // mm_interconnect_2:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                                      // hps_0:h2f_lw_WLAST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                      // mm_interconnect_2:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                       // hps_0:h2f_lw_AWID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                        // mm_interconnect_2:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                                     // mm_interconnect_2:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                     // hps_0:h2f_lw_AWSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                                    // hps_0:h2f_lw_AWVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                                     // mm_interconnect_2:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_2_dma_to_sdram_csr_readdata;                        // DMA_to_SDRAM:csr_readdata -> mm_interconnect_2:DMA_to_SDRAM_csr_readdata
	wire    [2:0] mm_interconnect_2_dma_to_sdram_csr_address;                         // mm_interconnect_2:DMA_to_SDRAM_csr_address -> DMA_to_SDRAM:csr_address
	wire          mm_interconnect_2_dma_to_sdram_csr_read;                            // mm_interconnect_2:DMA_to_SDRAM_csr_read -> DMA_to_SDRAM:csr_read
	wire    [3:0] mm_interconnect_2_dma_to_sdram_csr_byteenable;                      // mm_interconnect_2:DMA_to_SDRAM_csr_byteenable -> DMA_to_SDRAM:csr_byteenable
	wire          mm_interconnect_2_dma_to_sdram_csr_write;                           // mm_interconnect_2:DMA_to_SDRAM_csr_write -> DMA_to_SDRAM:csr_write
	wire   [31:0] mm_interconnect_2_dma_to_sdram_csr_writedata;                       // mm_interconnect_2:DMA_to_SDRAM_csr_writedata -> DMA_to_SDRAM:csr_writedata
	wire          mm_interconnect_2_dma_to_sdram_descriptor_slave_waitrequest;        // DMA_to_SDRAM:descriptor_slave_waitrequest -> mm_interconnect_2:DMA_to_SDRAM_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_2_dma_to_sdram_descriptor_slave_byteenable;         // mm_interconnect_2:DMA_to_SDRAM_descriptor_slave_byteenable -> DMA_to_SDRAM:descriptor_slave_byteenable
	wire          mm_interconnect_2_dma_to_sdram_descriptor_slave_write;              // mm_interconnect_2:DMA_to_SDRAM_descriptor_slave_write -> DMA_to_SDRAM:descriptor_slave_write
	wire  [127:0] mm_interconnect_2_dma_to_sdram_descriptor_slave_writedata;          // mm_interconnect_2:DMA_to_SDRAM_descriptor_slave_writedata -> DMA_to_SDRAM:descriptor_slave_writedata
	wire          pulsegenerator_cdc_m0_waitrequest;                                  // mm_interconnect_3:pulsegenerator_cdc_m0_waitrequest -> pulsegenerator_cdc:m0_waitrequest
	wire   [31:0] pulsegenerator_cdc_m0_readdata;                                     // mm_interconnect_3:pulsegenerator_cdc_m0_readdata -> pulsegenerator_cdc:m0_readdata
	wire          pulsegenerator_cdc_m0_debugaccess;                                  // pulsegenerator_cdc:m0_debugaccess -> mm_interconnect_3:pulsegenerator_cdc_m0_debugaccess
	wire    [3:0] pulsegenerator_cdc_m0_address;                                      // pulsegenerator_cdc:m0_address -> mm_interconnect_3:pulsegenerator_cdc_m0_address
	wire          pulsegenerator_cdc_m0_read;                                         // pulsegenerator_cdc:m0_read -> mm_interconnect_3:pulsegenerator_cdc_m0_read
	wire    [3:0] pulsegenerator_cdc_m0_byteenable;                                   // pulsegenerator_cdc:m0_byteenable -> mm_interconnect_3:pulsegenerator_cdc_m0_byteenable
	wire          pulsegenerator_cdc_m0_readdatavalid;                                // mm_interconnect_3:pulsegenerator_cdc_m0_readdatavalid -> pulsegenerator_cdc:m0_readdatavalid
	wire   [31:0] pulsegenerator_cdc_m0_writedata;                                    // pulsegenerator_cdc:m0_writedata -> mm_interconnect_3:pulsegenerator_cdc_m0_writedata
	wire          pulsegenerator_cdc_m0_write;                                        // pulsegenerator_cdc:m0_write -> mm_interconnect_3:pulsegenerator_cdc_m0_write
	wire    [0:0] pulsegenerator_cdc_m0_burstcount;                                   // pulsegenerator_cdc:m0_burstcount -> mm_interconnect_3:pulsegenerator_cdc_m0_burstcount
	wire    [3:0] mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awaddr;      // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_awaddr -> pulsegenerator:S_AXI_AWADDR
	wire    [1:0] mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_bresp;       // pulsegenerator:S_AXI_BRESP -> mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_bresp
	wire          mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_arready;     // pulsegenerator:S_AXI_ARREADY -> mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_arready
	wire   [31:0] mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rdata;       // pulsegenerator:S_AXI_RDATA -> mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_rdata
	wire    [3:0] mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wstrb;       // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_wstrb -> pulsegenerator:S_AXI_WSTRB
	wire          mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wready;      // pulsegenerator:S_AXI_WREADY -> mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_wready
	wire          mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awready;     // pulsegenerator:S_AXI_AWREADY -> mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_awready
	wire          mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rready;      // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_rready -> pulsegenerator:S_AXI_RREADY
	wire          mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_bready;      // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_bready -> pulsegenerator:S_AXI_BREADY
	wire          mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wvalid;      // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_wvalid -> pulsegenerator:S_AXI_WVALID
	wire    [3:0] mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_araddr;      // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_araddr -> pulsegenerator:S_AXI_ARADDR
	wire    [2:0] mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_arprot;      // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_arprot -> pulsegenerator:S_AXI_ARPROT
	wire    [1:0] mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rresp;       // pulsegenerator:S_AXI_RRESP -> mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_rresp
	wire    [2:0] mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awprot;      // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_awprot -> pulsegenerator:S_AXI_AWPROT
	wire   [31:0] mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wdata;       // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_wdata -> pulsegenerator:S_AXI_WDATA
	wire          mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_arvalid;     // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_arvalid -> pulsegenerator:S_AXI_ARVALID
	wire          mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_bvalid;      // pulsegenerator:S_AXI_BVALID -> mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_bvalid
	wire          mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awvalid;     // mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_awvalid -> pulsegenerator:S_AXI_AWVALID
	wire          mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rvalid;      // pulsegenerator:S_AXI_RVALID -> mm_interconnect_3:pulsegenerator_altera_axi4lite_slave_rvalid
	wire          ipsync_bridge_m0_waitrequest;                                       // mm_interconnect_4:ipsync_bridge_m0_waitrequest -> ipsync_bridge:m0_waitrequest
	wire   [31:0] ipsync_bridge_m0_readdata;                                          // mm_interconnect_4:ipsync_bridge_m0_readdata -> ipsync_bridge:m0_readdata
	wire          ipsync_bridge_m0_debugaccess;                                       // ipsync_bridge:m0_debugaccess -> mm_interconnect_4:ipsync_bridge_m0_debugaccess
	wire    [9:0] ipsync_bridge_m0_address;                                           // ipsync_bridge:m0_address -> mm_interconnect_4:ipsync_bridge_m0_address
	wire          ipsync_bridge_m0_read;                                              // ipsync_bridge:m0_read -> mm_interconnect_4:ipsync_bridge_m0_read
	wire    [3:0] ipsync_bridge_m0_byteenable;                                        // ipsync_bridge:m0_byteenable -> mm_interconnect_4:ipsync_bridge_m0_byteenable
	wire          ipsync_bridge_m0_readdatavalid;                                     // mm_interconnect_4:ipsync_bridge_m0_readdatavalid -> ipsync_bridge:m0_readdatavalid
	wire   [31:0] ipsync_bridge_m0_writedata;                                         // ipsync_bridge:m0_writedata -> mm_interconnect_4:ipsync_bridge_m0_writedata
	wire          ipsync_bridge_m0_write;                                             // ipsync_bridge:m0_write -> mm_interconnect_4:ipsync_bridge_m0_write
	wire    [0:0] ipsync_bridge_m0_burstcount;                                        // ipsync_bridge:m0_burstcount -> mm_interconnect_4:ipsync_bridge_m0_burstcount
	wire   [31:0] mm_interconnect_4_ip_sync_avalon_slave_readdata;                    // ip_sync:S_AVMM_RDATA -> mm_interconnect_4:ip_sync_avalon_slave_readdata
	wire          mm_interconnect_4_ip_sync_avalon_slave_waitrequest;                 // ip_sync:S_AVMM_WAITREQUEST -> mm_interconnect_4:ip_sync_avalon_slave_waitrequest
	wire    [7:0] mm_interconnect_4_ip_sync_avalon_slave_address;                     // mm_interconnect_4:ip_sync_avalon_slave_address -> ip_sync:S_AVMM_ADDR
	wire          mm_interconnect_4_ip_sync_avalon_slave_read;                        // mm_interconnect_4:ip_sync_avalon_slave_read -> ip_sync:S_AVMM_R
	wire    [3:0] mm_interconnect_4_ip_sync_avalon_slave_byteenable;                  // mm_interconnect_4:ip_sync_avalon_slave_byteenable -> ip_sync:S_AVMM_BYTEENABLE
	wire          mm_interconnect_4_ip_sync_avalon_slave_readdatavalid;               // ip_sync:S_AVMM_READATAVALID -> mm_interconnect_4:ip_sync_avalon_slave_readdatavalid
	wire          mm_interconnect_4_ip_sync_avalon_slave_write;                       // mm_interconnect_4:ip_sync_avalon_slave_write -> ip_sync:S_AVMM_W
	wire   [31:0] mm_interconnect_4_ip_sync_avalon_slave_writedata;                   // mm_interconnect_4:ip_sync_avalon_slave_writedata -> ip_sync:S_AVMM_WDATA
	wire    [0:0] mm_interconnect_4_ip_sync_avalon_slave_burstcount;                  // mm_interconnect_4:ip_sync_avalon_slave_burstcount -> ip_sync:S_AVMM_BURSTCOUNT
	wire          ipsync_to_aes_delay_m0_waitrequest;                                 // mm_interconnect_5:ipsync_to_aes_delay_m0_waitrequest -> ipsync_to_aes_delay:m0_waitrequest
	wire   [31:0] ipsync_to_aes_delay_m0_readdata;                                    // mm_interconnect_5:ipsync_to_aes_delay_m0_readdata -> ipsync_to_aes_delay:m0_readdata
	wire          ipsync_to_aes_delay_m0_debugaccess;                                 // ipsync_to_aes_delay:m0_debugaccess -> mm_interconnect_5:ipsync_to_aes_delay_m0_debugaccess
	wire    [9:0] ipsync_to_aes_delay_m0_address;                                     // ipsync_to_aes_delay:m0_address -> mm_interconnect_5:ipsync_to_aes_delay_m0_address
	wire          ipsync_to_aes_delay_m0_read;                                        // ipsync_to_aes_delay:m0_read -> mm_interconnect_5:ipsync_to_aes_delay_m0_read
	wire    [3:0] ipsync_to_aes_delay_m0_byteenable;                                  // ipsync_to_aes_delay:m0_byteenable -> mm_interconnect_5:ipsync_to_aes_delay_m0_byteenable
	wire          ipsync_to_aes_delay_m0_readdatavalid;                               // mm_interconnect_5:ipsync_to_aes_delay_m0_readdatavalid -> ipsync_to_aes_delay:m0_readdatavalid
	wire   [31:0] ipsync_to_aes_delay_m0_writedata;                                   // ipsync_to_aes_delay:m0_writedata -> mm_interconnect_5:ipsync_to_aes_delay_m0_writedata
	wire          ipsync_to_aes_delay_m0_write;                                       // ipsync_to_aes_delay:m0_write -> mm_interconnect_5:ipsync_to_aes_delay_m0_write
	wire    [0:0] ipsync_to_aes_delay_m0_burstcount;                                  // ipsync_to_aes_delay:m0_burstcount -> mm_interconnect_5:ipsync_to_aes_delay_m0_burstcount
	wire          mm_interconnect_5_aes_avalon_slave_0_1_chipselect;                  // mm_interconnect_5:aes_avalon_slave_0_1_chipselect -> aes:cs
	wire   [31:0] mm_interconnect_5_aes_avalon_slave_0_1_readdata;                    // aes:read_data -> mm_interconnect_5:aes_avalon_slave_0_1_readdata
	wire    [7:0] mm_interconnect_5_aes_avalon_slave_0_1_address;                     // mm_interconnect_5:aes_avalon_slave_0_1_address -> aes:address
	wire          mm_interconnect_5_aes_avalon_slave_0_1_write;                       // mm_interconnect_5:aes_avalon_slave_0_1_write -> aes:we
	wire   [31:0] mm_interconnect_5_aes_avalon_slave_0_1_writedata;                   // mm_interconnect_5:aes_avalon_slave_0_1_writedata -> aes:write_data
	wire          theta_pll_reconfig_cdc_m0_waitrequest;                              // mm_interconnect_6:theta_pll_reconfig_cdc_m0_waitrequest -> theta_pll_reconfig_cdc:m0_waitrequest
	wire   [31:0] theta_pll_reconfig_cdc_m0_readdata;                                 // mm_interconnect_6:theta_pll_reconfig_cdc_m0_readdata -> theta_pll_reconfig_cdc:m0_readdata
	wire          theta_pll_reconfig_cdc_m0_debugaccess;                              // theta_pll_reconfig_cdc:m0_debugaccess -> mm_interconnect_6:theta_pll_reconfig_cdc_m0_debugaccess
	wire    [7:0] theta_pll_reconfig_cdc_m0_address;                                  // theta_pll_reconfig_cdc:m0_address -> mm_interconnect_6:theta_pll_reconfig_cdc_m0_address
	wire          theta_pll_reconfig_cdc_m0_read;                                     // theta_pll_reconfig_cdc:m0_read -> mm_interconnect_6:theta_pll_reconfig_cdc_m0_read
	wire    [3:0] theta_pll_reconfig_cdc_m0_byteenable;                               // theta_pll_reconfig_cdc:m0_byteenable -> mm_interconnect_6:theta_pll_reconfig_cdc_m0_byteenable
	wire          theta_pll_reconfig_cdc_m0_readdatavalid;                            // mm_interconnect_6:theta_pll_reconfig_cdc_m0_readdatavalid -> theta_pll_reconfig_cdc:m0_readdatavalid
	wire   [31:0] theta_pll_reconfig_cdc_m0_writedata;                                // theta_pll_reconfig_cdc:m0_writedata -> mm_interconnect_6:theta_pll_reconfig_cdc_m0_writedata
	wire          theta_pll_reconfig_cdc_m0_write;                                    // theta_pll_reconfig_cdc:m0_write -> mm_interconnect_6:theta_pll_reconfig_cdc_m0_write
	wire    [0:0] theta_pll_reconfig_cdc_m0_burstcount;                               // theta_pll_reconfig_cdc:m0_burstcount -> mm_interconnect_6:theta_pll_reconfig_cdc_m0_burstcount
	wire   [31:0] mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_readdata;    // theta_pll_reconfig:mgmt_readdata -> mm_interconnect_6:theta_pll_reconfig_mgmt_avalon_slave_readdata
	wire          mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_waitrequest; // theta_pll_reconfig:mgmt_waitrequest -> mm_interconnect_6:theta_pll_reconfig_mgmt_avalon_slave_waitrequest
	wire    [5:0] mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_address;     // mm_interconnect_6:theta_pll_reconfig_mgmt_avalon_slave_address -> theta_pll_reconfig:mgmt_address
	wire          mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_read;        // mm_interconnect_6:theta_pll_reconfig_mgmt_avalon_slave_read -> theta_pll_reconfig:mgmt_read
	wire          mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_write;       // mm_interconnect_6:theta_pll_reconfig_mgmt_avalon_slave_write -> theta_pll_reconfig:mgmt_write
	wire   [31:0] mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_writedata;   // mm_interconnect_6:theta_pll_reconfig_mgmt_avalon_slave_writedata -> theta_pll_reconfig:mgmt_writedata
	wire          phi_pll_reconfig_cdc_m0_waitrequest;                                // mm_interconnect_7:phi_pll_reconfig_cdc_m0_waitrequest -> phi_pll_reconfig_cdc:m0_waitrequest
	wire   [31:0] phi_pll_reconfig_cdc_m0_readdata;                                   // mm_interconnect_7:phi_pll_reconfig_cdc_m0_readdata -> phi_pll_reconfig_cdc:m0_readdata
	wire          phi_pll_reconfig_cdc_m0_debugaccess;                                // phi_pll_reconfig_cdc:m0_debugaccess -> mm_interconnect_7:phi_pll_reconfig_cdc_m0_debugaccess
	wire    [7:0] phi_pll_reconfig_cdc_m0_address;                                    // phi_pll_reconfig_cdc:m0_address -> mm_interconnect_7:phi_pll_reconfig_cdc_m0_address
	wire          phi_pll_reconfig_cdc_m0_read;                                       // phi_pll_reconfig_cdc:m0_read -> mm_interconnect_7:phi_pll_reconfig_cdc_m0_read
	wire    [3:0] phi_pll_reconfig_cdc_m0_byteenable;                                 // phi_pll_reconfig_cdc:m0_byteenable -> mm_interconnect_7:phi_pll_reconfig_cdc_m0_byteenable
	wire          phi_pll_reconfig_cdc_m0_readdatavalid;                              // mm_interconnect_7:phi_pll_reconfig_cdc_m0_readdatavalid -> phi_pll_reconfig_cdc:m0_readdatavalid
	wire   [31:0] phi_pll_reconfig_cdc_m0_writedata;                                  // phi_pll_reconfig_cdc:m0_writedata -> mm_interconnect_7:phi_pll_reconfig_cdc_m0_writedata
	wire          phi_pll_reconfig_cdc_m0_write;                                      // phi_pll_reconfig_cdc:m0_write -> mm_interconnect_7:phi_pll_reconfig_cdc_m0_write
	wire    [0:0] phi_pll_reconfig_cdc_m0_burstcount;                                 // phi_pll_reconfig_cdc:m0_burstcount -> mm_interconnect_7:phi_pll_reconfig_cdc_m0_burstcount
	wire   [31:0] mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_readdata;      // phi_pll_reconfig:mgmt_readdata -> mm_interconnect_7:phi_pll_reconfig_mgmt_avalon_slave_readdata
	wire          mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_waitrequest;   // phi_pll_reconfig:mgmt_waitrequest -> mm_interconnect_7:phi_pll_reconfig_mgmt_avalon_slave_waitrequest
	wire    [5:0] mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_address;       // mm_interconnect_7:phi_pll_reconfig_mgmt_avalon_slave_address -> phi_pll_reconfig:mgmt_address
	wire          mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_read;          // mm_interconnect_7:phi_pll_reconfig_mgmt_avalon_slave_read -> phi_pll_reconfig:mgmt_read
	wire          mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_write;         // mm_interconnect_7:phi_pll_reconfig_mgmt_avalon_slave_write -> phi_pll_reconfig:mgmt_write
	wire   [31:0] mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_writedata;     // mm_interconnect_7:phi_pll_reconfig_mgmt_avalon_slave_writedata -> phi_pll_reconfig:mgmt_writedata
	wire          dma_to_sdram_mm_write_waitrequest;                                  // mm_interconnect_8:DMA_to_SDRAM_mm_write_waitrequest -> DMA_to_SDRAM:mm_write_waitrequest
	wire   [31:0] dma_to_sdram_mm_write_address;                                      // DMA_to_SDRAM:mm_write_address -> mm_interconnect_8:DMA_to_SDRAM_mm_write_address
	wire   [31:0] dma_to_sdram_mm_write_byteenable;                                   // DMA_to_SDRAM:mm_write_byteenable -> mm_interconnect_8:DMA_to_SDRAM_mm_write_byteenable
	wire          dma_to_sdram_mm_write_write;                                        // DMA_to_SDRAM:mm_write_write -> mm_interconnect_8:DMA_to_SDRAM_mm_write_write
	wire  [255:0] dma_to_sdram_mm_write_writedata;                                    // DMA_to_SDRAM:mm_write_writedata -> mm_interconnect_8:DMA_to_SDRAM_mm_write_writedata
	wire    [3:0] dma_to_sdram_mm_write_burstcount;                                   // DMA_to_SDRAM:mm_write_burstcount -> mm_interconnect_8:DMA_to_SDRAM_mm_write_burstcount
	wire          mm_interconnect_8_hps_0_f2h_sdram0_data_waitrequest;                // hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_8:hps_0_f2h_sdram0_data_waitrequest
	wire   [26:0] mm_interconnect_8_hps_0_f2h_sdram0_data_address;                    // mm_interconnect_8:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	wire   [31:0] mm_interconnect_8_hps_0_f2h_sdram0_data_byteenable;                 // mm_interconnect_8:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	wire          mm_interconnect_8_hps_0_f2h_sdram0_data_write;                      // mm_interconnect_8:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	wire  [255:0] mm_interconnect_8_hps_0_f2h_sdram0_data_writedata;                  // mm_interconnect_8:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	wire    [7:0] mm_interconnect_8_hps_0_f2h_sdram0_data_burstcount;                 // mm_interconnect_8:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	wire          irq_mapper_receiver0_irq;                                           // DMA_to_SDRAM:csr_irq_irq -> irq_mapper:receiver0_irq
	wire   [31:0] hps_0_f2h_irq0_irq;                                                 // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                                 // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [DMA_to_SDRAM:reset_n_reset_n, aes_reset_pio:reset_n, ipsync_bridge:s0_reset, mm_interconnect_1:theta_pll_reconfig_cdc_s0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:DMA_to_SDRAM_reset_n_reset_bridge_in_reset_reset, mm_interconnect_8:DMA_to_SDRAM_reset_n_reset_bridge_in_reset_reset, phi_locked:reset_n, phi_pll_reconfig_cdc:s0_reset, phi_pll_reset_pio:reset_n, tdc_reset_pio:reset_n, theta_locked:reset_n, theta_pll_reconfig_cdc:s0_reset, theta_pll_reset_pio:reset_n]
	wire          rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [aes:reset_n, ip_sync:reset, ipsync_bridge:m0_reset, ipsync_to_aes_delay:m0_reset, ipsync_to_aes_delay:s0_reset, mm_interconnect_0:ip_sync_reset_reset_bridge_in_reset_reset, mm_interconnect_4:ipsync_bridge_m0_reset_reset_bridge_in_reset_reset, mm_interconnect_5:ipsync_to_aes_delay_m0_reset_reset_bridge_in_reset_reset]
	wire          aes_reset_controller_reset_out_reset;                               // aes_reset_controller:reset_out -> rst_controller_001:reset_in2
	wire          rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> ip_sync_to_pulsegenerator_cdc:in_reset_n
	wire          rst_controller_003_reset_out_reset;                                 // rst_controller_003:reset_out -> ip_sync_to_pulsegenerator_cdc:out_reset_n
	wire          rst_controller_004_reset_out_reset;                                 // rst_controller_004:reset_out -> phi_clk:rst
	wire          phi_pll_reset_bridge_reset_out_reset;                               // phi_pll_reset_bridge:reset_out -> rst_controller_004:reset_in2
	wire          rst_controller_005_reset_out_reset;                                 // rst_controller_005:reset_out -> [mm_interconnect_6:theta_pll_reconfig_cdc_m0_reset_reset_bridge_in_reset_reset, mm_interconnect_7:phi_pll_reconfig_cdc_m0_reset_reset_bridge_in_reset_reset, phi_pll_reconfig:mgmt_reset, phi_pll_reconfig_cdc:m0_reset, theta_pll_reconfig:mgmt_reset, theta_pll_reconfig_cdc:m0_reset]
	wire          rst_controller_006_reset_out_reset;                                 // rst_controller_006:reset_out -> [mm_interconnect_3:pulsegenerator_cdc_m0_reset_reset_bridge_in_reset_reset, pulsegenerator:S_AXI_ARESETN, pulsegenerator_cdc:m0_reset]
	wire          reset_bridge_launch_reset_out_reset;                                // reset_bridge_launch:reset_out -> rst_controller_006:reset_in2
	wire          rst_controller_007_reset_out_reset;                                 // rst_controller_007:reset_out -> [mm_interconnect_1:pulsegenerator_cdc_s0_reset_reset_bridge_in_reset_reset, pulsegenerator_cdc:s0_reset, tdc_to_dma_dc_fifo:out_reset_n]
	wire          reset_bridge_shell_reset_out_reset;                                 // reset_bridge_shell:reset_out -> rst_controller_007:reset_in2
	wire          rst_controller_008_reset_out_reset;                                 // rst_controller_008:reset_out -> [tdc_0:reset, tdc_to_dma_dc_fifo:in_reset_n]
	wire          reset_bridge_capt_reset_out_reset;                                  // reset_bridge_capt:reset_out -> rst_controller_008:reset_in2
	wire          rst_controller_009_reset_out_reset;                                 // rst_controller_009:reset_out -> theta_clks:rst
	wire          theta_pll_reset_bridge_reset_out_reset;                             // theta_pll_reset_bridge:reset_out -> rst_controller_009:reset_in2
	wire          rst_controller_010_reset_out_reset;                                 // rst_controller_010:reset_out -> [mm_interconnect_1:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_8:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset]

	soc_system_DMA_to_SDRAM dma_to_sdram (
		.mm_write_address             (dma_to_sdram_mm_write_address),                               //         mm_write.address
		.mm_write_write               (dma_to_sdram_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (dma_to_sdram_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (dma_to_sdram_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (dma_to_sdram_mm_write_waitrequest),                           //                 .waitrequest
		.mm_write_burstcount          (dma_to_sdram_mm_write_burstcount),                            //                 .burstcount
		.clock_clk                    (shell_pll_outclk0_clk),                                       //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                             //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_2_dma_to_sdram_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_2_dma_to_sdram_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_2_dma_to_sdram_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_2_dma_to_sdram_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_2_dma_to_sdram_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_2_dma_to_sdram_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_2_dma_to_sdram_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_2_dma_to_sdram_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_2_dma_to_sdram_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_2_dma_to_sdram_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_receiver0_irq),                                    //          csr_irq.irq
		.st_sink_data                 (tdc_to_dma_dc_fifo_out_data),                                 //          st_sink.data
		.st_sink_valid                (tdc_to_dma_dc_fifo_out_valid),                                //                 .valid
		.st_sink_ready                (tdc_to_dma_dc_fifo_out_ready)                                 //                 .ready
	);

	aes aes (
		.clk        (shell_pll_outclk1_clk),                             //            clock.clk
		.reset_n    (~rst_controller_001_reset_out_reset),               //            reset.reset_n
		.cs         (mm_interconnect_5_aes_avalon_slave_0_1_chipselect), // avalon_slave_0_1.chipselect
		.we         (mm_interconnect_5_aes_avalon_slave_0_1_write),      //                 .write
		.address    (mm_interconnect_5_aes_avalon_slave_0_1_address),    //                 .address
		.write_data (mm_interconnect_5_aes_avalon_slave_0_1_writedata),  //                 .writedata
		.read_data  (mm_interconnect_5_aes_avalon_slave_0_1_readdata)    //                 .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) aes_reset_controller (
		.reset_in0      (aes_reset_in_reset),                   // reset_in0.reset
		.clk            (shell_pll_outclk1_clk),                //       clk.clk
		.reset_out      (aes_reset_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_in1      (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	soc_system_aes_reset_pio aes_reset_pio (
		.clk        (shell_pll_outclk0_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_1_aes_reset_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_aes_reset_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_aes_reset_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_aes_reset_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_aes_reset_pio_s1_readdata),   //                    .readdata
		.out_port   (aes_reset_out_export)                           // external_connection.export
	);

	soc_system_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.mem_a                  (memory_mem_a),                                        //            memory.mem_a
		.mem_ba                 (memory_mem_ba),                                       //                  .mem_ba
		.mem_ck                 (memory_mem_ck),                                       //                  .mem_ck
		.mem_ck_n               (memory_mem_ck_n),                                     //                  .mem_ck_n
		.mem_cke                (memory_mem_cke),                                      //                  .mem_cke
		.mem_cs_n               (memory_mem_cs_n),                                     //                  .mem_cs_n
		.mem_ras_n              (memory_mem_ras_n),                                    //                  .mem_ras_n
		.mem_cas_n              (memory_mem_cas_n),                                    //                  .mem_cas_n
		.mem_we_n               (memory_mem_we_n),                                     //                  .mem_we_n
		.mem_reset_n            (memory_mem_reset_n),                                  //                  .mem_reset_n
		.mem_dq                 (memory_mem_dq),                                       //                  .mem_dq
		.mem_dqs                (memory_mem_dqs),                                      //                  .mem_dqs
		.mem_dqs_n              (memory_mem_dqs_n),                                    //                  .mem_dqs_n
		.mem_odt                (memory_mem_odt),                                      //                  .mem_odt
		.mem_dm                 (memory_mem_dm),                                       //                  .mem_dm
		.oct_rzqin              (memory_oct_rzqin),                                    //                  .oct_rzqin
		.h2f_rst_n              (hps_0_h2f_reset_reset),                               //         h2f_reset.reset_n
		.f2h_sdram0_clk         (shell_pll_outclk0_clk),                               //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS     (mm_interconnect_8_hps_0_f2h_sdram0_data_address),     //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT  (mm_interconnect_8_hps_0_f2h_sdram0_data_burstcount),  //                  .burstcount
		.f2h_sdram0_WAITREQUEST (mm_interconnect_8_hps_0_f2h_sdram0_data_waitrequest), //                  .waitrequest
		.f2h_sdram0_WRITEDATA   (mm_interconnect_8_hps_0_f2h_sdram0_data_writedata),   //                  .writedata
		.f2h_sdram0_BYTEENABLE  (mm_interconnect_8_hps_0_f2h_sdram0_data_byteenable),  //                  .byteenable
		.f2h_sdram0_WRITE       (mm_interconnect_8_hps_0_f2h_sdram0_data_write),       //                  .write
		.h2f_axi_clk            (shell_pll_outclk0_clk),                               //     h2f_axi_clock.clk
		.h2f_AWID               (hps_0_h2f_axi_master_awid),                           //    h2f_axi_master.awid
		.h2f_AWADDR             (hps_0_h2f_axi_master_awaddr),                         //                  .awaddr
		.h2f_AWLEN              (hps_0_h2f_axi_master_awlen),                          //                  .awlen
		.h2f_AWSIZE             (hps_0_h2f_axi_master_awsize),                         //                  .awsize
		.h2f_AWBURST            (hps_0_h2f_axi_master_awburst),                        //                  .awburst
		.h2f_AWLOCK             (hps_0_h2f_axi_master_awlock),                         //                  .awlock
		.h2f_AWCACHE            (hps_0_h2f_axi_master_awcache),                        //                  .awcache
		.h2f_AWPROT             (hps_0_h2f_axi_master_awprot),                         //                  .awprot
		.h2f_AWVALID            (hps_0_h2f_axi_master_awvalid),                        //                  .awvalid
		.h2f_AWREADY            (hps_0_h2f_axi_master_awready),                        //                  .awready
		.h2f_WID                (hps_0_h2f_axi_master_wid),                            //                  .wid
		.h2f_WDATA              (hps_0_h2f_axi_master_wdata),                          //                  .wdata
		.h2f_WSTRB              (hps_0_h2f_axi_master_wstrb),                          //                  .wstrb
		.h2f_WLAST              (hps_0_h2f_axi_master_wlast),                          //                  .wlast
		.h2f_WVALID             (hps_0_h2f_axi_master_wvalid),                         //                  .wvalid
		.h2f_WREADY             (hps_0_h2f_axi_master_wready),                         //                  .wready
		.h2f_BID                (hps_0_h2f_axi_master_bid),                            //                  .bid
		.h2f_BRESP              (hps_0_h2f_axi_master_bresp),                          //                  .bresp
		.h2f_BVALID             (hps_0_h2f_axi_master_bvalid),                         //                  .bvalid
		.h2f_BREADY             (hps_0_h2f_axi_master_bready),                         //                  .bready
		.h2f_ARID               (hps_0_h2f_axi_master_arid),                           //                  .arid
		.h2f_ARADDR             (hps_0_h2f_axi_master_araddr),                         //                  .araddr
		.h2f_ARLEN              (hps_0_h2f_axi_master_arlen),                          //                  .arlen
		.h2f_ARSIZE             (hps_0_h2f_axi_master_arsize),                         //                  .arsize
		.h2f_ARBURST            (hps_0_h2f_axi_master_arburst),                        //                  .arburst
		.h2f_ARLOCK             (hps_0_h2f_axi_master_arlock),                         //                  .arlock
		.h2f_ARCACHE            (hps_0_h2f_axi_master_arcache),                        //                  .arcache
		.h2f_ARPROT             (hps_0_h2f_axi_master_arprot),                         //                  .arprot
		.h2f_ARVALID            (hps_0_h2f_axi_master_arvalid),                        //                  .arvalid
		.h2f_ARREADY            (hps_0_h2f_axi_master_arready),                        //                  .arready
		.h2f_RID                (hps_0_h2f_axi_master_rid),                            //                  .rid
		.h2f_RDATA              (hps_0_h2f_axi_master_rdata),                          //                  .rdata
		.h2f_RRESP              (hps_0_h2f_axi_master_rresp),                          //                  .rresp
		.h2f_RLAST              (hps_0_h2f_axi_master_rlast),                          //                  .rlast
		.h2f_RVALID             (hps_0_h2f_axi_master_rvalid),                         //                  .rvalid
		.h2f_RREADY             (hps_0_h2f_axi_master_rready),                         //                  .rready
		.h2f_lw_axi_clk         (shell_pll_outclk0_clk),                               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID            (hps_0_h2f_lw_axi_master_awid),                        // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR          (hps_0_h2f_lw_axi_master_awaddr),                      //                  .awaddr
		.h2f_lw_AWLEN           (hps_0_h2f_lw_axi_master_awlen),                       //                  .awlen
		.h2f_lw_AWSIZE          (hps_0_h2f_lw_axi_master_awsize),                      //                  .awsize
		.h2f_lw_AWBURST         (hps_0_h2f_lw_axi_master_awburst),                     //                  .awburst
		.h2f_lw_AWLOCK          (hps_0_h2f_lw_axi_master_awlock),                      //                  .awlock
		.h2f_lw_AWCACHE         (hps_0_h2f_lw_axi_master_awcache),                     //                  .awcache
		.h2f_lw_AWPROT          (hps_0_h2f_lw_axi_master_awprot),                      //                  .awprot
		.h2f_lw_AWVALID         (hps_0_h2f_lw_axi_master_awvalid),                     //                  .awvalid
		.h2f_lw_AWREADY         (hps_0_h2f_lw_axi_master_awready),                     //                  .awready
		.h2f_lw_WID             (hps_0_h2f_lw_axi_master_wid),                         //                  .wid
		.h2f_lw_WDATA           (hps_0_h2f_lw_axi_master_wdata),                       //                  .wdata
		.h2f_lw_WSTRB           (hps_0_h2f_lw_axi_master_wstrb),                       //                  .wstrb
		.h2f_lw_WLAST           (hps_0_h2f_lw_axi_master_wlast),                       //                  .wlast
		.h2f_lw_WVALID          (hps_0_h2f_lw_axi_master_wvalid),                      //                  .wvalid
		.h2f_lw_WREADY          (hps_0_h2f_lw_axi_master_wready),                      //                  .wready
		.h2f_lw_BID             (hps_0_h2f_lw_axi_master_bid),                         //                  .bid
		.h2f_lw_BRESP           (hps_0_h2f_lw_axi_master_bresp),                       //                  .bresp
		.h2f_lw_BVALID          (hps_0_h2f_lw_axi_master_bvalid),                      //                  .bvalid
		.h2f_lw_BREADY          (hps_0_h2f_lw_axi_master_bready),                      //                  .bready
		.h2f_lw_ARID            (hps_0_h2f_lw_axi_master_arid),                        //                  .arid
		.h2f_lw_ARADDR          (hps_0_h2f_lw_axi_master_araddr),                      //                  .araddr
		.h2f_lw_ARLEN           (hps_0_h2f_lw_axi_master_arlen),                       //                  .arlen
		.h2f_lw_ARSIZE          (hps_0_h2f_lw_axi_master_arsize),                      //                  .arsize
		.h2f_lw_ARBURST         (hps_0_h2f_lw_axi_master_arburst),                     //                  .arburst
		.h2f_lw_ARLOCK          (hps_0_h2f_lw_axi_master_arlock),                      //                  .arlock
		.h2f_lw_ARCACHE         (hps_0_h2f_lw_axi_master_arcache),                     //                  .arcache
		.h2f_lw_ARPROT          (hps_0_h2f_lw_axi_master_arprot),                      //                  .arprot
		.h2f_lw_ARVALID         (hps_0_h2f_lw_axi_master_arvalid),                     //                  .arvalid
		.h2f_lw_ARREADY         (hps_0_h2f_lw_axi_master_arready),                     //                  .arready
		.h2f_lw_RID             (hps_0_h2f_lw_axi_master_rid),                         //                  .rid
		.h2f_lw_RDATA           (hps_0_h2f_lw_axi_master_rdata),                       //                  .rdata
		.h2f_lw_RRESP           (hps_0_h2f_lw_axi_master_rresp),                       //                  .rresp
		.h2f_lw_RLAST           (hps_0_h2f_lw_axi_master_rlast),                       //                  .rlast
		.h2f_lw_RVALID          (hps_0_h2f_lw_axi_master_rvalid),                      //                  .rvalid
		.h2f_lw_RREADY          (hps_0_h2f_lw_axi_master_rready),                      //                  .rready
		.f2h_irq_p0             (hps_0_f2h_irq0_irq),                                  //          f2h_irq0.irq
		.f2h_irq_p1             (hps_0_f2h_irq1_irq)                                   //          f2h_irq1.irq
	);

	ip_sync #(
		.ADDR_TRIGGER (9'b000001000),
		.DATA_TRIGGER (34'b0000000000000000000000000000000010)
	) ip_sync (
		.reset               (rst_controller_001_reset_out_reset),                   //                   reset.reset
		.clk                 (shell_pll_outclk1_clk),                                //                   clock.clk
		.M_AVMM_ADDR         (ip_sync_avalon_master_address),                        //           avalon_master.address
		.M_AVMM_RDATA        (ip_sync_avalon_master_readdata),                       //                        .readdata
		.M_AVMM_W            (ip_sync_avalon_master_write),                          //                        .write
		.M_AVMM_WDATA        (ip_sync_avalon_master_writedata),                      //                        .writedata
		.M_AVMM_WAITREQUEST  (ip_sync_avalon_master_waitrequest),                    //                        .waitrequest
		.M_AVMM_BURSTCOUNT   (ip_sync_avalon_master_burstcount),                     //                        .burstcount
		.M_AVMM_BYTEENABLE   (ip_sync_avalon_master_byteenable),                     //                        .byteenable
		.M_AVMM_READATAVALID (ip_sync_avalon_master_readdatavalid),                  //                        .readdatavalid
		.M_AVMM_R            (ip_sync_avalon_master_read),                           //                        .read
		.S_AVMM_ADDR         (mm_interconnect_4_ip_sync_avalon_slave_address),       //            avalon_slave.address
		.S_AVMM_RDATA        (mm_interconnect_4_ip_sync_avalon_slave_readdata),      //                        .readdata
		.S_AVMM_W            (mm_interconnect_4_ip_sync_avalon_slave_write),         //                        .write
		.S_AVMM_WDATA        (mm_interconnect_4_ip_sync_avalon_slave_writedata),     //                        .writedata
		.S_AVMM_WAITREQUEST  (mm_interconnect_4_ip_sync_avalon_slave_waitrequest),   //                        .waitrequest
		.S_AVMM_R            (mm_interconnect_4_ip_sync_avalon_slave_read),          //                        .read
		.S_AVMM_READATAVALID (mm_interconnect_4_ip_sync_avalon_slave_readdatavalid), //                        .readdatavalid
		.S_AVMM_BURSTCOUNT   (mm_interconnect_4_ip_sync_avalon_slave_burstcount),    //                        .burstcount
		.S_AVMM_BYTEENABLE   (mm_interconnect_4_ip_sync_avalon_slave_byteenable),    //                        .byteenable
		.M_AVST_DATA         (ip_sync_avalon_streaming_source_data),                 // avalon_streaming_source.data
		.M_AVST_READY        (ip_sync_avalon_streaming_source_ready),                //                        .ready
		.M_AVST_VALID        (ip_sync_avalon_streaming_source_valid)                 //                        .valid
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (16),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (0),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (8),
		.RD_SYNC_DEPTH      (8)
	) ip_sync_to_pulsegenerator_cdc (
		.in_clk            (shell_pll_outclk1_clk),                   //        in_clk.clk
		.in_reset_n        (~rst_controller_002_reset_out_reset),     //  in_clk_reset.reset_n
		.out_clk           (theta_clks_outclk0_clk),                  //       out_clk.clk
		.out_reset_n       (~rst_controller_003_reset_out_reset),     // out_clk_reset.reset_n
		.in_data           (ip_sync_avalon_streaming_source_data),    //            in.data
		.in_valid          (ip_sync_avalon_streaming_source_valid),   //              .valid
		.in_ready          (ip_sync_avalon_streaming_source_ready),   //              .ready
		.out_data          (ip_sync_to_pulsegenerator_cdc_out_data),  //           out.data
		.out_valid         (ip_sync_to_pulsegenerator_cdc_out_valid), //              .valid
		.out_ready         (ip_sync_to_pulsegenerator_cdc_out_ready), //              .ready
		.in_csr_address    (1'b0),                                    //   (terminated)
		.in_csr_read       (1'b0),                                    //   (terminated)
		.in_csr_write      (1'b0),                                    //   (terminated)
		.in_csr_readdata   (),                                        //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000),    //   (terminated)
		.out_csr_address   (1'b0),                                    //   (terminated)
		.out_csr_read      (1'b0),                                    //   (terminated)
		.out_csr_write     (1'b0),                                    //   (terminated)
		.out_csr_readdata  (),                                        //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000),    //   (terminated)
		.in_startofpacket  (1'b0),                                    //   (terminated)
		.in_endofpacket    (1'b0),                                    //   (terminated)
		.out_startofpacket (),                                        //   (terminated)
		.out_endofpacket   (),                                        //   (terminated)
		.in_empty          (1'b0),                                    //   (terminated)
		.out_empty         (),                                        //   (terminated)
		.in_error          (1'b0),                                    //   (terminated)
		.out_error         (),                                        //   (terminated)
		.in_channel        (1'b0),                                    //   (terminated)
		.out_channel       (),                                        //   (terminated)
		.space_avail_data  ()                                         //   (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (8),
		.MASTER_SYNC_DEPTH   (8),
		.SLAVE_SYNC_DEPTH    (8)
	) ipsync_bridge (
		.m0_clk           (shell_pll_outclk1_clk),                            //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),               // m0_reset.reset
		.s0_clk           (shell_pll_outclk0_clk),                            //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                   // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_1_ipsync_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_1_ipsync_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_1_ipsync_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_1_ipsync_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_1_ipsync_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_1_ipsync_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_1_ipsync_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_1_ipsync_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_1_ipsync_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_1_ipsync_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (ipsync_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (ipsync_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (ipsync_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (ipsync_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (ipsync_bridge_m0_writedata),                       //         .writedata
		.m0_address       (ipsync_bridge_m0_address),                         //         .address
		.m0_write         (ipsync_bridge_m0_write),                           //         .write
		.m0_read          (ipsync_bridge_m0_read),                            //         .read
		.m0_byteenable    (ipsync_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (ipsync_bridge_m0_debugaccess)                      //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (8),
		.MASTER_SYNC_DEPTH   (16),
		.SLAVE_SYNC_DEPTH    (16)
	) ipsync_to_aes_delay (
		.m0_clk           (shell_pll_outclk1_clk),                                  //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                     // m0_reset.reset
		.s0_clk           (shell_pll_outclk1_clk),                                  //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                     // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_ipsync_to_aes_delay_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_ipsync_to_aes_delay_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_ipsync_to_aes_delay_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_ipsync_to_aes_delay_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_ipsync_to_aes_delay_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_ipsync_to_aes_delay_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_ipsync_to_aes_delay_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_ipsync_to_aes_delay_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_ipsync_to_aes_delay_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_ipsync_to_aes_delay_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (ipsync_to_aes_delay_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (ipsync_to_aes_delay_m0_readdata),                        //         .readdata
		.m0_readdatavalid (ipsync_to_aes_delay_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (ipsync_to_aes_delay_m0_burstcount),                      //         .burstcount
		.m0_writedata     (ipsync_to_aes_delay_m0_writedata),                       //         .writedata
		.m0_address       (ipsync_to_aes_delay_m0_address),                         //         .address
		.m0_write         (ipsync_to_aes_delay_m0_write),                           //         .write
		.m0_read          (ipsync_to_aes_delay_m0_read),                            //         .read
		.m0_byteenable    (ipsync_to_aes_delay_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (ipsync_to_aes_delay_m0_debugaccess)                      //         .debugaccess
	);

	soc_system_phi_clk phi_clk (
		.refclk            (clk_clk),                                          //            refclk.clk
		.rst               (rst_controller_004_reset_out_reset),               //             reset.reset
		.outclk_0          (),                                                 //           outclk0.clk
		.locked            (locked_phi_out_export),                            //            locked.export
		.cascade_out       (phi_clk_cascade_out_export),                       //       cascade_out.export
		.reconfig_to_pll   (phi_pll_reconfig_reconfig_to_pll_reconfig_to_pll), //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (phi_clk_reconfig_from_pll_reconfig_from_pll)       // reconfig_from_pll.reconfig_from_pll
	);

	soc_system_phi_locked phi_locked (
		.clk      (shell_pll_outclk0_clk),                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_phi_locked_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_phi_locked_s1_readdata), //                    .readdata
		.in_port  (locked_phi_in_export)                      // external_connection.export
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) phi_pll_reconfig (
		.mgmt_clk          (clk_clk),                                                          //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_005_reset_out_reset),                               //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (phi_pll_reconfig_reconfig_to_pll_reconfig_to_pll),                 //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (phi_clk_reconfig_from_pll_reconfig_from_pll),                      // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                           //       (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (8),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (8),
		.MASTER_SYNC_DEPTH   (8),
		.SLAVE_SYNC_DEPTH    (8)
	) phi_pll_reconfig_cdc (
		.m0_clk           (clk_clk),                                                 //   m0_clk.clk
		.m0_reset         (rst_controller_005_reset_out_reset),                      // m0_reset.reset
		.s0_clk           (shell_pll_outclk0_clk),                                   //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                          // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_1_phi_pll_reconfig_cdc_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_1_phi_pll_reconfig_cdc_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_1_phi_pll_reconfig_cdc_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_1_phi_pll_reconfig_cdc_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_1_phi_pll_reconfig_cdc_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_1_phi_pll_reconfig_cdc_s0_address),       //         .address
		.s0_write         (mm_interconnect_1_phi_pll_reconfig_cdc_s0_write),         //         .write
		.s0_read          (mm_interconnect_1_phi_pll_reconfig_cdc_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_1_phi_pll_reconfig_cdc_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_1_phi_pll_reconfig_cdc_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (phi_pll_reconfig_cdc_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (phi_pll_reconfig_cdc_m0_readdata),                        //         .readdata
		.m0_readdatavalid (phi_pll_reconfig_cdc_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (phi_pll_reconfig_cdc_m0_burstcount),                      //         .burstcount
		.m0_writedata     (phi_pll_reconfig_cdc_m0_writedata),                       //         .writedata
		.m0_address       (phi_pll_reconfig_cdc_m0_address),                         //         .address
		.m0_write         (phi_pll_reconfig_cdc_m0_write),                           //         .write
		.m0_read          (phi_pll_reconfig_cdc_m0_read),                            //         .read
		.m0_byteenable    (phi_pll_reconfig_cdc_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (phi_pll_reconfig_cdc_m0_debugaccess)                      //         .debugaccess
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) phi_pll_reset_bridge (
		.reset_in0      (reset_phi_in_reset),                   // reset_in0.reset
		.clk            (clk_clk),                              //       clk.clk
		.reset_out      (phi_pll_reset_bridge_reset_out_reset), // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_in1      (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	soc_system_aes_reset_pio phi_pll_reset_pio (
		.clk        (shell_pll_outclk0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_1_phi_pll_reset_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_phi_pll_reset_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_phi_pll_reset_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_phi_pll_reset_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_phi_pll_reset_pio_s1_readdata),   //                    .readdata
		.out_port   (reset_phi_out_export)                               // external_connection.export
	);

	pulsegenerator #(
		.C_SELECT_BIT    (4'b0001),
		.PIPELINE_OUTPUT (4)
	) pulsegenerator (
		.S_AXI_ACLK    (theta_clks_outclk0_clk),                                         //             axi_s_clock.clk
		.S_AXI_ARESETN (~rst_controller_006_reset_out_reset),                            //            axi_s_resetn.reset_n
		.S_AXI_ARADDR  (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_araddr),  //   altera_axi4lite_slave.araddr
		.S_AXI_ARREADY (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_arready), //                        .arready
		.S_AXI_ARVALID (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_arvalid), //                        .arvalid
		.S_AXI_AWADDR  (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awaddr),  //                        .awaddr
		.S_AXI_AWREADY (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awready), //                        .awready
		.S_AXI_AWVALID (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awvalid), //                        .awvalid
		.S_AXI_BREADY  (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_bready),  //                        .bready
		.S_AXI_BRESP   (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_bresp),   //                        .bresp
		.S_AXI_BVALID  (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_bvalid),  //                        .bvalid
		.S_AXI_RDATA   (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rdata),   //                        .rdata
		.S_AXI_RREADY  (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rready),  //                        .rready
		.S_AXI_RRESP   (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rresp),   //                        .rresp
		.S_AXI_RVALID  (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rvalid),  //                        .rvalid
		.S_AXI_WDATA   (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wdata),   //                        .wdata
		.S_AXI_WREADY  (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wready),  //                        .wready
		.S_AXI_WSTRB   (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wstrb),   //                        .wstrb
		.S_AXI_WVALID  (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wvalid),  //                        .wvalid
		.S_AXI_ARPROT  (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_arprot),  //                        .arprot
		.S_AXI_AWPROT  (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awprot),  //                        .awprot
		.M_AVST_DATA   (pulsegenerator_avalon_streaming_source_data),                    // avalon_streaming_source.data
		.M_AVST_VALID  (pulsegenerator_avalon_streaming_source_valid),                   //                        .valid
		.M_AVST_READY  (pulsegenerator_avalon_streaming_source_ready),                   //                        .ready
		.S_AVST_VALID  (ip_sync_to_pulsegenerator_cdc_out_valid),                        //   avalon_streaming_sink.valid
		.S_AVST_DATA   (ip_sync_to_pulsegenerator_cdc_out_data),                         //                        .data
		.S_AVST_READY  (ip_sync_to_pulsegenerator_cdc_out_ready)                         //                        .ready
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (4),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (8),
		.MASTER_SYNC_DEPTH   (8),
		.SLAVE_SYNC_DEPTH    (8)
	) pulsegenerator_cdc (
		.m0_clk           (theta_clks_outclk0_clk),                                //   m0_clk.clk
		.m0_reset         (rst_controller_006_reset_out_reset),                    // m0_reset.reset
		.s0_clk           (shell_pll_outclk0_clk),                                 //   s0_clk.clk
		.s0_reset         (rst_controller_007_reset_out_reset),                    // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_1_pulsegenerator_cdc_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_1_pulsegenerator_cdc_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_1_pulsegenerator_cdc_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_1_pulsegenerator_cdc_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_1_pulsegenerator_cdc_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_1_pulsegenerator_cdc_s0_address),       //         .address
		.s0_write         (mm_interconnect_1_pulsegenerator_cdc_s0_write),         //         .write
		.s0_read          (mm_interconnect_1_pulsegenerator_cdc_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_1_pulsegenerator_cdc_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_1_pulsegenerator_cdc_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (pulsegenerator_cdc_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (pulsegenerator_cdc_m0_readdata),                        //         .readdata
		.m0_readdatavalid (pulsegenerator_cdc_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (pulsegenerator_cdc_m0_burstcount),                      //         .burstcount
		.m0_writedata     (pulsegenerator_cdc_m0_writedata),                       //         .writedata
		.m0_address       (pulsegenerator_cdc_m0_address),                         //         .address
		.m0_write         (pulsegenerator_cdc_m0_write),                           //         .write
		.m0_read          (pulsegenerator_cdc_m0_read),                            //         .read
		.m0_byteenable    (pulsegenerator_cdc_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (pulsegenerator_cdc_m0_debugaccess)                      //         .debugaccess
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_bridge_capt (
		.reset_in0      (reset_bridge_tdc_reset_out_reset),  // reset_in0.reset
		.clk            (theta_clks_outclk1_clk),            //       clk.clk
		.reset_out      (reset_bridge_capt_reset_out_reset), // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_in1      (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_bridge_launch (
		.reset_in0      (reset_bridge_tdc_reset_out_reset),    // reset_in0.reset
		.clk            (theta_clks_outclk0_clk),              //       clk.clk
		.reset_out      (reset_bridge_launch_reset_out_reset), // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_bridge_shell (
		.reset_in0      (reset_bridge_tdc_reset_out_reset),   // reset_in0.reset
		.clk            (shell_pll_outclk0_clk),              //       clk.clk
		.reset_out      (reset_bridge_shell_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_bridge_tdc (
		.reset_in0      (tdc_reset_in_reset),               // reset_in0.reset
		.clk            (shell_pll_outclk0_clk),            //       clk.clk
		.reset_out      (reset_bridge_tdc_reset_out_reset), // reset_out.reset
		.reset_req      (),                                 // (terminated)
		.reset_req_in0  (1'b0),                             // (terminated)
		.reset_in1      (1'b0),                             // (terminated)
		.reset_req_in1  (1'b0),                             // (terminated)
		.reset_in2      (1'b0),                             // (terminated)
		.reset_req_in2  (1'b0),                             // (terminated)
		.reset_in3      (1'b0),                             // (terminated)
		.reset_req_in3  (1'b0),                             // (terminated)
		.reset_in4      (1'b0),                             // (terminated)
		.reset_req_in4  (1'b0),                             // (terminated)
		.reset_in5      (1'b0),                             // (terminated)
		.reset_req_in5  (1'b0),                             // (terminated)
		.reset_in6      (1'b0),                             // (terminated)
		.reset_req_in6  (1'b0),                             // (terminated)
		.reset_in7      (1'b0),                             // (terminated)
		.reset_req_in7  (1'b0),                             // (terminated)
		.reset_in8      (1'b0),                             // (terminated)
		.reset_req_in8  (1'b0),                             // (terminated)
		.reset_in9      (1'b0),                             // (terminated)
		.reset_req_in9  (1'b0),                             // (terminated)
		.reset_in10     (1'b0),                             // (terminated)
		.reset_req_in10 (1'b0),                             // (terminated)
		.reset_in11     (1'b0),                             // (terminated)
		.reset_req_in11 (1'b0),                             // (terminated)
		.reset_in12     (1'b0),                             // (terminated)
		.reset_req_in12 (1'b0),                             // (terminated)
		.reset_in13     (1'b0),                             // (terminated)
		.reset_req_in13 (1'b0),                             // (terminated)
		.reset_in14     (1'b0),                             // (terminated)
		.reset_req_in14 (1'b0),                             // (terminated)
		.reset_in15     (1'b0),                             // (terminated)
		.reset_req_in15 (1'b0)                              // (terminated)
	);

	soc_system_shell_pll shell_pll (
		.refclk   (clk_clk),                //  refclk.clk
		.rst      (~hps_0_h2f_reset_reset), //   reset.reset
		.outclk_0 (shell_pll_outclk0_clk),  // outclk0.clk
		.outclk_1 (shell_pll_outclk1_clk),  // outclk1.clk
		.locked   ()                        // (terminated)
	);

	tdc_top #(
		.C_OUT_WIDTH  (128),
		.C_SYNC_DEPTH (4),
		.TECHNOLOGY   ("28nm"),
		.REVERSE      (1)
	) tdc_0 (
		.reset        (rst_controller_008_reset_out_reset),           //                   reset.reset
		.clk_capt     (theta_clks_outclk1_clk),                       //                clk_capt.clk
		.clk_launch   (theta_clks_outclk0_clk),                       //              clk_launch.clk
		.S_AVST_DATA  (pulsegenerator_avalon_streaming_source_data),  //   avalon_streaming_sink.data
		.S_AVST_VALID (pulsegenerator_avalon_streaming_source_valid), //                        .valid
		.S_AVST_READY (pulsegenerator_avalon_streaming_source_ready), //                        .ready
		.M_AVST_DATA  (tdc_0_avalon_streaming_source_data),           // avalon_streaming_source.data
		.M_AVST_VALID (tdc_0_avalon_streaming_source_valid),          //                        .valid
		.M_AVST_READY (tdc_0_avalon_streaming_source_ready)           //                        .ready
	);

	soc_system_aes_reset_pio tdc_reset_pio (
		.clk        (shell_pll_outclk0_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_1_tdc_reset_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_tdc_reset_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_tdc_reset_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_tdc_reset_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_tdc_reset_pio_s1_readdata),   //                    .readdata
		.out_port   (tdc_reset_out_export)                           // external_connection.export
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (32),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (16),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (0),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (8),
		.RD_SYNC_DEPTH      (8)
	) tdc_to_dma_dc_fifo (
		.in_clk            (theta_clks_outclk1_clk),               //        in_clk.clk
		.in_reset_n        (~rst_controller_008_reset_out_reset),  //  in_clk_reset.reset_n
		.out_clk           (shell_pll_outclk0_clk),                //       out_clk.clk
		.out_reset_n       (~rst_controller_007_reset_out_reset),  // out_clk_reset.reset_n
		.in_data           (tdc_0_avalon_streaming_source_data),   //            in.data
		.in_valid          (tdc_0_avalon_streaming_source_valid),  //              .valid
		.in_ready          (tdc_0_avalon_streaming_source_ready),  //              .ready
		.out_data          (tdc_to_dma_dc_fifo_out_data),          //           out.data
		.out_valid         (tdc_to_dma_dc_fifo_out_valid),         //              .valid
		.out_ready         (tdc_to_dma_dc_fifo_out_ready),         //              .ready
		.in_csr_address    (1'b0),                                 //   (terminated)
		.in_csr_read       (1'b0),                                 //   (terminated)
		.in_csr_write      (1'b0),                                 //   (terminated)
		.in_csr_readdata   (),                                     //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000), //   (terminated)
		.out_csr_address   (1'b0),                                 //   (terminated)
		.out_csr_read      (1'b0),                                 //   (terminated)
		.out_csr_write     (1'b0),                                 //   (terminated)
		.out_csr_readdata  (),                                     //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000), //   (terminated)
		.in_startofpacket  (1'b0),                                 //   (terminated)
		.in_endofpacket    (1'b0),                                 //   (terminated)
		.out_startofpacket (),                                     //   (terminated)
		.out_endofpacket   (),                                     //   (terminated)
		.in_empty          (5'b00000),                             //   (terminated)
		.out_empty         (),                                     //   (terminated)
		.in_error          (1'b0),                                 //   (terminated)
		.out_error         (),                                     //   (terminated)
		.in_channel        (1'b0),                                 //   (terminated)
		.out_channel       (),                                     //   (terminated)
		.space_avail_data  ()                                      //   (terminated)
	);

	soc_system_theta_clks theta_clks (
		.refclk            (theta_clks_refclk_clk),                              //            refclk.clk
		.rst               (rst_controller_009_reset_out_reset),                 //             reset.reset
		.outclk_0          (theta_clks_outclk0_clk),                             //           outclk0.clk
		.outclk_1          (theta_clks_outclk1_clk),                             //           outclk1.clk
		.locked            (locked_theta_out_export),                            //            locked.export
		.adjpllin          (phi_clk_cascade_out_export),                         //          adjpllin.export
		.reconfig_to_pll   (theta_pll_reconfig_reconfig_to_pll_reconfig_to_pll), //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (theta_clks_reconfig_from_pll_reconfig_from_pll)      // reconfig_from_pll.reconfig_from_pll
	);

	soc_system_phi_locked theta_locked (
		.clk      (shell_pll_outclk0_clk),                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_theta_locked_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_theta_locked_s1_readdata), //                    .readdata
		.in_port  (locked_theta_in_export)                      // external_connection.export
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) theta_pll_reconfig (
		.mgmt_clk          (clk_clk),                                                            //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_005_reset_out_reset),                                 //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (theta_pll_reconfig_reconfig_to_pll_reconfig_to_pll),                 //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (theta_clks_reconfig_from_pll_reconfig_from_pll),                     // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                             //       (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (8),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (8),
		.MASTER_SYNC_DEPTH   (8),
		.SLAVE_SYNC_DEPTH    (8)
	) theta_pll_reconfig_cdc (
		.m0_clk           (clk_clk),                                                   //   m0_clk.clk
		.m0_reset         (rst_controller_005_reset_out_reset),                        // m0_reset.reset
		.s0_clk           (shell_pll_outclk0_clk),                                     //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                            // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_1_theta_pll_reconfig_cdc_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_1_theta_pll_reconfig_cdc_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_1_theta_pll_reconfig_cdc_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_1_theta_pll_reconfig_cdc_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_1_theta_pll_reconfig_cdc_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_1_theta_pll_reconfig_cdc_s0_address),       //         .address
		.s0_write         (mm_interconnect_1_theta_pll_reconfig_cdc_s0_write),         //         .write
		.s0_read          (mm_interconnect_1_theta_pll_reconfig_cdc_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_1_theta_pll_reconfig_cdc_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_1_theta_pll_reconfig_cdc_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (theta_pll_reconfig_cdc_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (theta_pll_reconfig_cdc_m0_readdata),                        //         .readdata
		.m0_readdatavalid (theta_pll_reconfig_cdc_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (theta_pll_reconfig_cdc_m0_burstcount),                      //         .burstcount
		.m0_writedata     (theta_pll_reconfig_cdc_m0_writedata),                       //         .writedata
		.m0_address       (theta_pll_reconfig_cdc_m0_address),                         //         .address
		.m0_write         (theta_pll_reconfig_cdc_m0_write),                           //         .write
		.m0_read          (theta_pll_reconfig_cdc_m0_read),                            //         .read
		.m0_byteenable    (theta_pll_reconfig_cdc_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (theta_pll_reconfig_cdc_m0_debugaccess)                      //         .debugaccess
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) theta_pll_reset_bridge (
		.reset_in0      (reset_theta_in_reset),                   // reset_in0.reset
		.clk            (shell_pll_outclk0_clk),                  //       clk.clk
		.reset_out      (theta_pll_reset_bridge_reset_out_reset), // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	soc_system_aes_reset_pio theta_pll_reset_pio (
		.clk        (shell_pll_outclk0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (mm_interconnect_1_theta_pll_reset_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_theta_pll_reset_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_theta_pll_reset_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_theta_pll_reset_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_theta_pll_reset_pio_s1_readdata),   //                    .readdata
		.out_port   (reset_theta_out_export)                               // external_connection.export
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.shell_pll_outclk1_clk                     (shell_pll_outclk1_clk),                                  //                   shell_pll_outclk1.clk
		.ip_sync_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                     // ip_sync_reset_reset_bridge_in_reset.reset
		.ip_sync_avalon_master_address             (ip_sync_avalon_master_address),                          //               ip_sync_avalon_master.address
		.ip_sync_avalon_master_waitrequest         (ip_sync_avalon_master_waitrequest),                      //                                    .waitrequest
		.ip_sync_avalon_master_burstcount          (ip_sync_avalon_master_burstcount),                       //                                    .burstcount
		.ip_sync_avalon_master_byteenable          (ip_sync_avalon_master_byteenable),                       //                                    .byteenable
		.ip_sync_avalon_master_read                (ip_sync_avalon_master_read),                             //                                    .read
		.ip_sync_avalon_master_readdata            (ip_sync_avalon_master_readdata),                         //                                    .readdata
		.ip_sync_avalon_master_readdatavalid       (ip_sync_avalon_master_readdatavalid),                    //                                    .readdatavalid
		.ip_sync_avalon_master_write               (ip_sync_avalon_master_write),                            //                                    .write
		.ip_sync_avalon_master_writedata           (ip_sync_avalon_master_writedata),                        //                                    .writedata
		.ipsync_to_aes_delay_s0_address            (mm_interconnect_0_ipsync_to_aes_delay_s0_address),       //              ipsync_to_aes_delay_s0.address
		.ipsync_to_aes_delay_s0_write              (mm_interconnect_0_ipsync_to_aes_delay_s0_write),         //                                    .write
		.ipsync_to_aes_delay_s0_read               (mm_interconnect_0_ipsync_to_aes_delay_s0_read),          //                                    .read
		.ipsync_to_aes_delay_s0_readdata           (mm_interconnect_0_ipsync_to_aes_delay_s0_readdata),      //                                    .readdata
		.ipsync_to_aes_delay_s0_writedata          (mm_interconnect_0_ipsync_to_aes_delay_s0_writedata),     //                                    .writedata
		.ipsync_to_aes_delay_s0_burstcount         (mm_interconnect_0_ipsync_to_aes_delay_s0_burstcount),    //                                    .burstcount
		.ipsync_to_aes_delay_s0_byteenable         (mm_interconnect_0_ipsync_to_aes_delay_s0_byteenable),    //                                    .byteenable
		.ipsync_to_aes_delay_s0_readdatavalid      (mm_interconnect_0_ipsync_to_aes_delay_s0_readdatavalid), //                                    .readdatavalid
		.ipsync_to_aes_delay_s0_waitrequest        (mm_interconnect_0_ipsync_to_aes_delay_s0_waitrequest),   //                                    .waitrequest
		.ipsync_to_aes_delay_s0_debugaccess        (mm_interconnect_0_ipsync_to_aes_delay_s0_debugaccess)    //                                    .debugaccess
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                 //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                               //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                               //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                              //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                               //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                              //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                               //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                              //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                              //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                  //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                               //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                               //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                  //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                               //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                               //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                 //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                               //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                               //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                              //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                               //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                              //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                               //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                              //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                              //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                  //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                               //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                               //                                                           .rready
		.shell_pll_outclk0_clk                                            (shell_pll_outclk0_clk),                                     //                                          shell_pll_outclk0.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_010_reset_out_reset),                        // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.pulsegenerator_cdc_s0_reset_reset_bridge_in_reset_reset          (rst_controller_007_reset_out_reset),                        //          pulsegenerator_cdc_s0_reset_reset_bridge_in_reset.reset
		.theta_pll_reconfig_cdc_s0_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                            //      theta_pll_reconfig_cdc_s0_reset_reset_bridge_in_reset.reset
		.aes_reset_pio_s1_address                                         (mm_interconnect_1_aes_reset_pio_s1_address),                //                                           aes_reset_pio_s1.address
		.aes_reset_pio_s1_write                                           (mm_interconnect_1_aes_reset_pio_s1_write),                  //                                                           .write
		.aes_reset_pio_s1_readdata                                        (mm_interconnect_1_aes_reset_pio_s1_readdata),               //                                                           .readdata
		.aes_reset_pio_s1_writedata                                       (mm_interconnect_1_aes_reset_pio_s1_writedata),              //                                                           .writedata
		.aes_reset_pio_s1_chipselect                                      (mm_interconnect_1_aes_reset_pio_s1_chipselect),             //                                                           .chipselect
		.ipsync_bridge_s0_address                                         (mm_interconnect_1_ipsync_bridge_s0_address),                //                                           ipsync_bridge_s0.address
		.ipsync_bridge_s0_write                                           (mm_interconnect_1_ipsync_bridge_s0_write),                  //                                                           .write
		.ipsync_bridge_s0_read                                            (mm_interconnect_1_ipsync_bridge_s0_read),                   //                                                           .read
		.ipsync_bridge_s0_readdata                                        (mm_interconnect_1_ipsync_bridge_s0_readdata),               //                                                           .readdata
		.ipsync_bridge_s0_writedata                                       (mm_interconnect_1_ipsync_bridge_s0_writedata),              //                                                           .writedata
		.ipsync_bridge_s0_burstcount                                      (mm_interconnect_1_ipsync_bridge_s0_burstcount),             //                                                           .burstcount
		.ipsync_bridge_s0_byteenable                                      (mm_interconnect_1_ipsync_bridge_s0_byteenable),             //                                                           .byteenable
		.ipsync_bridge_s0_readdatavalid                                   (mm_interconnect_1_ipsync_bridge_s0_readdatavalid),          //                                                           .readdatavalid
		.ipsync_bridge_s0_waitrequest                                     (mm_interconnect_1_ipsync_bridge_s0_waitrequest),            //                                                           .waitrequest
		.ipsync_bridge_s0_debugaccess                                     (mm_interconnect_1_ipsync_bridge_s0_debugaccess),            //                                                           .debugaccess
		.phi_locked_s1_address                                            (mm_interconnect_1_phi_locked_s1_address),                   //                                              phi_locked_s1.address
		.phi_locked_s1_readdata                                           (mm_interconnect_1_phi_locked_s1_readdata),                  //                                                           .readdata
		.phi_pll_reconfig_cdc_s0_address                                  (mm_interconnect_1_phi_pll_reconfig_cdc_s0_address),         //                                    phi_pll_reconfig_cdc_s0.address
		.phi_pll_reconfig_cdc_s0_write                                    (mm_interconnect_1_phi_pll_reconfig_cdc_s0_write),           //                                                           .write
		.phi_pll_reconfig_cdc_s0_read                                     (mm_interconnect_1_phi_pll_reconfig_cdc_s0_read),            //                                                           .read
		.phi_pll_reconfig_cdc_s0_readdata                                 (mm_interconnect_1_phi_pll_reconfig_cdc_s0_readdata),        //                                                           .readdata
		.phi_pll_reconfig_cdc_s0_writedata                                (mm_interconnect_1_phi_pll_reconfig_cdc_s0_writedata),       //                                                           .writedata
		.phi_pll_reconfig_cdc_s0_burstcount                               (mm_interconnect_1_phi_pll_reconfig_cdc_s0_burstcount),      //                                                           .burstcount
		.phi_pll_reconfig_cdc_s0_byteenable                               (mm_interconnect_1_phi_pll_reconfig_cdc_s0_byteenable),      //                                                           .byteenable
		.phi_pll_reconfig_cdc_s0_readdatavalid                            (mm_interconnect_1_phi_pll_reconfig_cdc_s0_readdatavalid),   //                                                           .readdatavalid
		.phi_pll_reconfig_cdc_s0_waitrequest                              (mm_interconnect_1_phi_pll_reconfig_cdc_s0_waitrequest),     //                                                           .waitrequest
		.phi_pll_reconfig_cdc_s0_debugaccess                              (mm_interconnect_1_phi_pll_reconfig_cdc_s0_debugaccess),     //                                                           .debugaccess
		.phi_pll_reset_pio_s1_address                                     (mm_interconnect_1_phi_pll_reset_pio_s1_address),            //                                       phi_pll_reset_pio_s1.address
		.phi_pll_reset_pio_s1_write                                       (mm_interconnect_1_phi_pll_reset_pio_s1_write),              //                                                           .write
		.phi_pll_reset_pio_s1_readdata                                    (mm_interconnect_1_phi_pll_reset_pio_s1_readdata),           //                                                           .readdata
		.phi_pll_reset_pio_s1_writedata                                   (mm_interconnect_1_phi_pll_reset_pio_s1_writedata),          //                                                           .writedata
		.phi_pll_reset_pio_s1_chipselect                                  (mm_interconnect_1_phi_pll_reset_pio_s1_chipselect),         //                                                           .chipselect
		.pulsegenerator_cdc_s0_address                                    (mm_interconnect_1_pulsegenerator_cdc_s0_address),           //                                      pulsegenerator_cdc_s0.address
		.pulsegenerator_cdc_s0_write                                      (mm_interconnect_1_pulsegenerator_cdc_s0_write),             //                                                           .write
		.pulsegenerator_cdc_s0_read                                       (mm_interconnect_1_pulsegenerator_cdc_s0_read),              //                                                           .read
		.pulsegenerator_cdc_s0_readdata                                   (mm_interconnect_1_pulsegenerator_cdc_s0_readdata),          //                                                           .readdata
		.pulsegenerator_cdc_s0_writedata                                  (mm_interconnect_1_pulsegenerator_cdc_s0_writedata),         //                                                           .writedata
		.pulsegenerator_cdc_s0_burstcount                                 (mm_interconnect_1_pulsegenerator_cdc_s0_burstcount),        //                                                           .burstcount
		.pulsegenerator_cdc_s0_byteenable                                 (mm_interconnect_1_pulsegenerator_cdc_s0_byteenable),        //                                                           .byteenable
		.pulsegenerator_cdc_s0_readdatavalid                              (mm_interconnect_1_pulsegenerator_cdc_s0_readdatavalid),     //                                                           .readdatavalid
		.pulsegenerator_cdc_s0_waitrequest                                (mm_interconnect_1_pulsegenerator_cdc_s0_waitrequest),       //                                                           .waitrequest
		.pulsegenerator_cdc_s0_debugaccess                                (mm_interconnect_1_pulsegenerator_cdc_s0_debugaccess),       //                                                           .debugaccess
		.tdc_reset_pio_s1_address                                         (mm_interconnect_1_tdc_reset_pio_s1_address),                //                                           tdc_reset_pio_s1.address
		.tdc_reset_pio_s1_write                                           (mm_interconnect_1_tdc_reset_pio_s1_write),                  //                                                           .write
		.tdc_reset_pio_s1_readdata                                        (mm_interconnect_1_tdc_reset_pio_s1_readdata),               //                                                           .readdata
		.tdc_reset_pio_s1_writedata                                       (mm_interconnect_1_tdc_reset_pio_s1_writedata),              //                                                           .writedata
		.tdc_reset_pio_s1_chipselect                                      (mm_interconnect_1_tdc_reset_pio_s1_chipselect),             //                                                           .chipselect
		.theta_locked_s1_address                                          (mm_interconnect_1_theta_locked_s1_address),                 //                                            theta_locked_s1.address
		.theta_locked_s1_readdata                                         (mm_interconnect_1_theta_locked_s1_readdata),                //                                                           .readdata
		.theta_pll_reconfig_cdc_s0_address                                (mm_interconnect_1_theta_pll_reconfig_cdc_s0_address),       //                                  theta_pll_reconfig_cdc_s0.address
		.theta_pll_reconfig_cdc_s0_write                                  (mm_interconnect_1_theta_pll_reconfig_cdc_s0_write),         //                                                           .write
		.theta_pll_reconfig_cdc_s0_read                                   (mm_interconnect_1_theta_pll_reconfig_cdc_s0_read),          //                                                           .read
		.theta_pll_reconfig_cdc_s0_readdata                               (mm_interconnect_1_theta_pll_reconfig_cdc_s0_readdata),      //                                                           .readdata
		.theta_pll_reconfig_cdc_s0_writedata                              (mm_interconnect_1_theta_pll_reconfig_cdc_s0_writedata),     //                                                           .writedata
		.theta_pll_reconfig_cdc_s0_burstcount                             (mm_interconnect_1_theta_pll_reconfig_cdc_s0_burstcount),    //                                                           .burstcount
		.theta_pll_reconfig_cdc_s0_byteenable                             (mm_interconnect_1_theta_pll_reconfig_cdc_s0_byteenable),    //                                                           .byteenable
		.theta_pll_reconfig_cdc_s0_readdatavalid                          (mm_interconnect_1_theta_pll_reconfig_cdc_s0_readdatavalid), //                                                           .readdatavalid
		.theta_pll_reconfig_cdc_s0_waitrequest                            (mm_interconnect_1_theta_pll_reconfig_cdc_s0_waitrequest),   //                                                           .waitrequest
		.theta_pll_reconfig_cdc_s0_debugaccess                            (mm_interconnect_1_theta_pll_reconfig_cdc_s0_debugaccess),   //                                                           .debugaccess
		.theta_pll_reset_pio_s1_address                                   (mm_interconnect_1_theta_pll_reset_pio_s1_address),          //                                     theta_pll_reset_pio_s1.address
		.theta_pll_reset_pio_s1_write                                     (mm_interconnect_1_theta_pll_reset_pio_s1_write),            //                                                           .write
		.theta_pll_reset_pio_s1_readdata                                  (mm_interconnect_1_theta_pll_reset_pio_s1_readdata),         //                                                           .readdata
		.theta_pll_reset_pio_s1_writedata                                 (mm_interconnect_1_theta_pll_reset_pio_s1_writedata),        //                                                           .writedata
		.theta_pll_reset_pio_s1_chipselect                                (mm_interconnect_1_theta_pll_reset_pio_s1_chipselect)        //                                                           .chipselect
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                              //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                               //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                              //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                             //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                              //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                             //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                              //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                             //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                             //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                 //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                               //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                               //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                               //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                              //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                              //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                 //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                               //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                              //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                              //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                              //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                               //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                              //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                             //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                              //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                             //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                              //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                             //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                             //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                 //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                               //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                               //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                               //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                              //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                              //                                                              .rready
		.shell_pll_outclk0_clk                                               (shell_pll_outclk0_clk),                                       //                                             shell_pll_outclk0.clk
		.DMA_to_SDRAM_reset_n_reset_bridge_in_reset_reset                    (rst_controller_reset_out_reset),                              //                    DMA_to_SDRAM_reset_n_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_010_reset_out_reset),                          // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.DMA_to_SDRAM_csr_address                                            (mm_interconnect_2_dma_to_sdram_csr_address),                  //                                              DMA_to_SDRAM_csr.address
		.DMA_to_SDRAM_csr_write                                              (mm_interconnect_2_dma_to_sdram_csr_write),                    //                                                              .write
		.DMA_to_SDRAM_csr_read                                               (mm_interconnect_2_dma_to_sdram_csr_read),                     //                                                              .read
		.DMA_to_SDRAM_csr_readdata                                           (mm_interconnect_2_dma_to_sdram_csr_readdata),                 //                                                              .readdata
		.DMA_to_SDRAM_csr_writedata                                          (mm_interconnect_2_dma_to_sdram_csr_writedata),                //                                                              .writedata
		.DMA_to_SDRAM_csr_byteenable                                         (mm_interconnect_2_dma_to_sdram_csr_byteenable),               //                                                              .byteenable
		.DMA_to_SDRAM_descriptor_slave_write                                 (mm_interconnect_2_dma_to_sdram_descriptor_slave_write),       //                                 DMA_to_SDRAM_descriptor_slave.write
		.DMA_to_SDRAM_descriptor_slave_writedata                             (mm_interconnect_2_dma_to_sdram_descriptor_slave_writedata),   //                                                              .writedata
		.DMA_to_SDRAM_descriptor_slave_byteenable                            (mm_interconnect_2_dma_to_sdram_descriptor_slave_byteenable),  //                                                              .byteenable
		.DMA_to_SDRAM_descriptor_slave_waitrequest                           (mm_interconnect_2_dma_to_sdram_descriptor_slave_waitrequest)  //                                                              .waitrequest
	);

	soc_system_mm_interconnect_3 mm_interconnect_3 (
		.pulsegenerator_altera_axi4lite_slave_awaddr             (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awaddr),  //              pulsegenerator_altera_axi4lite_slave.awaddr
		.pulsegenerator_altera_axi4lite_slave_awprot             (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awprot),  //                                                  .awprot
		.pulsegenerator_altera_axi4lite_slave_awvalid            (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awvalid), //                                                  .awvalid
		.pulsegenerator_altera_axi4lite_slave_awready            (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_awready), //                                                  .awready
		.pulsegenerator_altera_axi4lite_slave_wdata              (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wdata),   //                                                  .wdata
		.pulsegenerator_altera_axi4lite_slave_wstrb              (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wstrb),   //                                                  .wstrb
		.pulsegenerator_altera_axi4lite_slave_wvalid             (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wvalid),  //                                                  .wvalid
		.pulsegenerator_altera_axi4lite_slave_wready             (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_wready),  //                                                  .wready
		.pulsegenerator_altera_axi4lite_slave_bresp              (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_bresp),   //                                                  .bresp
		.pulsegenerator_altera_axi4lite_slave_bvalid             (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_bvalid),  //                                                  .bvalid
		.pulsegenerator_altera_axi4lite_slave_bready             (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_bready),  //                                                  .bready
		.pulsegenerator_altera_axi4lite_slave_araddr             (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_araddr),  //                                                  .araddr
		.pulsegenerator_altera_axi4lite_slave_arprot             (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_arprot),  //                                                  .arprot
		.pulsegenerator_altera_axi4lite_slave_arvalid            (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_arvalid), //                                                  .arvalid
		.pulsegenerator_altera_axi4lite_slave_arready            (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_arready), //                                                  .arready
		.pulsegenerator_altera_axi4lite_slave_rdata              (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rdata),   //                                                  .rdata
		.pulsegenerator_altera_axi4lite_slave_rresp              (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rresp),   //                                                  .rresp
		.pulsegenerator_altera_axi4lite_slave_rvalid             (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rvalid),  //                                                  .rvalid
		.pulsegenerator_altera_axi4lite_slave_rready             (mm_interconnect_3_pulsegenerator_altera_axi4lite_slave_rready),  //                                                  .rready
		.theta_clks_outclk0_clk                                  (theta_clks_outclk0_clk),                                         //                                theta_clks_outclk0.clk
		.pulsegenerator_cdc_m0_reset_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),                             // pulsegenerator_cdc_m0_reset_reset_bridge_in_reset.reset
		.pulsegenerator_cdc_m0_address                           (pulsegenerator_cdc_m0_address),                                  //                             pulsegenerator_cdc_m0.address
		.pulsegenerator_cdc_m0_waitrequest                       (pulsegenerator_cdc_m0_waitrequest),                              //                                                  .waitrequest
		.pulsegenerator_cdc_m0_burstcount                        (pulsegenerator_cdc_m0_burstcount),                               //                                                  .burstcount
		.pulsegenerator_cdc_m0_byteenable                        (pulsegenerator_cdc_m0_byteenable),                               //                                                  .byteenable
		.pulsegenerator_cdc_m0_read                              (pulsegenerator_cdc_m0_read),                                     //                                                  .read
		.pulsegenerator_cdc_m0_readdata                          (pulsegenerator_cdc_m0_readdata),                                 //                                                  .readdata
		.pulsegenerator_cdc_m0_readdatavalid                     (pulsegenerator_cdc_m0_readdatavalid),                            //                                                  .readdatavalid
		.pulsegenerator_cdc_m0_write                             (pulsegenerator_cdc_m0_write),                                    //                                                  .write
		.pulsegenerator_cdc_m0_writedata                         (pulsegenerator_cdc_m0_writedata),                                //                                                  .writedata
		.pulsegenerator_cdc_m0_debugaccess                       (pulsegenerator_cdc_m0_debugaccess)                               //                                                  .debugaccess
	);

	soc_system_mm_interconnect_4 mm_interconnect_4 (
		.shell_pll_outclk1_clk                              (shell_pll_outclk1_clk),                                //                            shell_pll_outclk1.clk
		.ipsync_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                   // ipsync_bridge_m0_reset_reset_bridge_in_reset.reset
		.ipsync_bridge_m0_address                           (ipsync_bridge_m0_address),                             //                             ipsync_bridge_m0.address
		.ipsync_bridge_m0_waitrequest                       (ipsync_bridge_m0_waitrequest),                         //                                             .waitrequest
		.ipsync_bridge_m0_burstcount                        (ipsync_bridge_m0_burstcount),                          //                                             .burstcount
		.ipsync_bridge_m0_byteenable                        (ipsync_bridge_m0_byteenable),                          //                                             .byteenable
		.ipsync_bridge_m0_read                              (ipsync_bridge_m0_read),                                //                                             .read
		.ipsync_bridge_m0_readdata                          (ipsync_bridge_m0_readdata),                            //                                             .readdata
		.ipsync_bridge_m0_readdatavalid                     (ipsync_bridge_m0_readdatavalid),                       //                                             .readdatavalid
		.ipsync_bridge_m0_write                             (ipsync_bridge_m0_write),                               //                                             .write
		.ipsync_bridge_m0_writedata                         (ipsync_bridge_m0_writedata),                           //                                             .writedata
		.ipsync_bridge_m0_debugaccess                       (ipsync_bridge_m0_debugaccess),                         //                                             .debugaccess
		.ip_sync_avalon_slave_address                       (mm_interconnect_4_ip_sync_avalon_slave_address),       //                         ip_sync_avalon_slave.address
		.ip_sync_avalon_slave_write                         (mm_interconnect_4_ip_sync_avalon_slave_write),         //                                             .write
		.ip_sync_avalon_slave_read                          (mm_interconnect_4_ip_sync_avalon_slave_read),          //                                             .read
		.ip_sync_avalon_slave_readdata                      (mm_interconnect_4_ip_sync_avalon_slave_readdata),      //                                             .readdata
		.ip_sync_avalon_slave_writedata                     (mm_interconnect_4_ip_sync_avalon_slave_writedata),     //                                             .writedata
		.ip_sync_avalon_slave_burstcount                    (mm_interconnect_4_ip_sync_avalon_slave_burstcount),    //                                             .burstcount
		.ip_sync_avalon_slave_byteenable                    (mm_interconnect_4_ip_sync_avalon_slave_byteenable),    //                                             .byteenable
		.ip_sync_avalon_slave_readdatavalid                 (mm_interconnect_4_ip_sync_avalon_slave_readdatavalid), //                                             .readdatavalid
		.ip_sync_avalon_slave_waitrequest                   (mm_interconnect_4_ip_sync_avalon_slave_waitrequest)    //                                             .waitrequest
	);

	soc_system_mm_interconnect_5 mm_interconnect_5 (
		.shell_pll_outclk1_clk                                    (shell_pll_outclk1_clk),                             //                                  shell_pll_outclk1.clk
		.ipsync_to_aes_delay_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                // ipsync_to_aes_delay_m0_reset_reset_bridge_in_reset.reset
		.ipsync_to_aes_delay_m0_address                           (ipsync_to_aes_delay_m0_address),                    //                             ipsync_to_aes_delay_m0.address
		.ipsync_to_aes_delay_m0_waitrequest                       (ipsync_to_aes_delay_m0_waitrequest),                //                                                   .waitrequest
		.ipsync_to_aes_delay_m0_burstcount                        (ipsync_to_aes_delay_m0_burstcount),                 //                                                   .burstcount
		.ipsync_to_aes_delay_m0_byteenable                        (ipsync_to_aes_delay_m0_byteenable),                 //                                                   .byteenable
		.ipsync_to_aes_delay_m0_read                              (ipsync_to_aes_delay_m0_read),                       //                                                   .read
		.ipsync_to_aes_delay_m0_readdata                          (ipsync_to_aes_delay_m0_readdata),                   //                                                   .readdata
		.ipsync_to_aes_delay_m0_readdatavalid                     (ipsync_to_aes_delay_m0_readdatavalid),              //                                                   .readdatavalid
		.ipsync_to_aes_delay_m0_write                             (ipsync_to_aes_delay_m0_write),                      //                                                   .write
		.ipsync_to_aes_delay_m0_writedata                         (ipsync_to_aes_delay_m0_writedata),                  //                                                   .writedata
		.ipsync_to_aes_delay_m0_debugaccess                       (ipsync_to_aes_delay_m0_debugaccess),                //                                                   .debugaccess
		.aes_avalon_slave_0_1_address                             (mm_interconnect_5_aes_avalon_slave_0_1_address),    //                               aes_avalon_slave_0_1.address
		.aes_avalon_slave_0_1_write                               (mm_interconnect_5_aes_avalon_slave_0_1_write),      //                                                   .write
		.aes_avalon_slave_0_1_readdata                            (mm_interconnect_5_aes_avalon_slave_0_1_readdata),   //                                                   .readdata
		.aes_avalon_slave_0_1_writedata                           (mm_interconnect_5_aes_avalon_slave_0_1_writedata),  //                                                   .writedata
		.aes_avalon_slave_0_1_chipselect                          (mm_interconnect_5_aes_avalon_slave_0_1_chipselect)  //                                                   .chipselect
	);

	soc_system_mm_interconnect_6 mm_interconnect_6 (
		.input_clk_clk_clk                                           (clk_clk),                                                            //                                         input_clk_clk.clk
		.theta_pll_reconfig_cdc_m0_reset_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),                                 // theta_pll_reconfig_cdc_m0_reset_reset_bridge_in_reset.reset
		.theta_pll_reconfig_cdc_m0_address                           (theta_pll_reconfig_cdc_m0_address),                                  //                             theta_pll_reconfig_cdc_m0.address
		.theta_pll_reconfig_cdc_m0_waitrequest                       (theta_pll_reconfig_cdc_m0_waitrequest),                              //                                                      .waitrequest
		.theta_pll_reconfig_cdc_m0_burstcount                        (theta_pll_reconfig_cdc_m0_burstcount),                               //                                                      .burstcount
		.theta_pll_reconfig_cdc_m0_byteenable                        (theta_pll_reconfig_cdc_m0_byteenable),                               //                                                      .byteenable
		.theta_pll_reconfig_cdc_m0_read                              (theta_pll_reconfig_cdc_m0_read),                                     //                                                      .read
		.theta_pll_reconfig_cdc_m0_readdata                          (theta_pll_reconfig_cdc_m0_readdata),                                 //                                                      .readdata
		.theta_pll_reconfig_cdc_m0_readdatavalid                     (theta_pll_reconfig_cdc_m0_readdatavalid),                            //                                                      .readdatavalid
		.theta_pll_reconfig_cdc_m0_write                             (theta_pll_reconfig_cdc_m0_write),                                    //                                                      .write
		.theta_pll_reconfig_cdc_m0_writedata                         (theta_pll_reconfig_cdc_m0_writedata),                                //                                                      .writedata
		.theta_pll_reconfig_cdc_m0_debugaccess                       (theta_pll_reconfig_cdc_m0_debugaccess),                              //                                                      .debugaccess
		.theta_pll_reconfig_mgmt_avalon_slave_address                (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_address),     //                  theta_pll_reconfig_mgmt_avalon_slave.address
		.theta_pll_reconfig_mgmt_avalon_slave_write                  (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_write),       //                                                      .write
		.theta_pll_reconfig_mgmt_avalon_slave_read                   (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_read),        //                                                      .read
		.theta_pll_reconfig_mgmt_avalon_slave_readdata               (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_readdata),    //                                                      .readdata
		.theta_pll_reconfig_mgmt_avalon_slave_writedata              (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_writedata),   //                                                      .writedata
		.theta_pll_reconfig_mgmt_avalon_slave_waitrequest            (mm_interconnect_6_theta_pll_reconfig_mgmt_avalon_slave_waitrequest)  //                                                      .waitrequest
	);

	soc_system_mm_interconnect_7 mm_interconnect_7 (
		.input_clk_clk_clk                                         (clk_clk),                                                          //                                       input_clk_clk.clk
		.phi_pll_reconfig_cdc_m0_reset_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),                               // phi_pll_reconfig_cdc_m0_reset_reset_bridge_in_reset.reset
		.phi_pll_reconfig_cdc_m0_address                           (phi_pll_reconfig_cdc_m0_address),                                  //                             phi_pll_reconfig_cdc_m0.address
		.phi_pll_reconfig_cdc_m0_waitrequest                       (phi_pll_reconfig_cdc_m0_waitrequest),                              //                                                    .waitrequest
		.phi_pll_reconfig_cdc_m0_burstcount                        (phi_pll_reconfig_cdc_m0_burstcount),                               //                                                    .burstcount
		.phi_pll_reconfig_cdc_m0_byteenable                        (phi_pll_reconfig_cdc_m0_byteenable),                               //                                                    .byteenable
		.phi_pll_reconfig_cdc_m0_read                              (phi_pll_reconfig_cdc_m0_read),                                     //                                                    .read
		.phi_pll_reconfig_cdc_m0_readdata                          (phi_pll_reconfig_cdc_m0_readdata),                                 //                                                    .readdata
		.phi_pll_reconfig_cdc_m0_readdatavalid                     (phi_pll_reconfig_cdc_m0_readdatavalid),                            //                                                    .readdatavalid
		.phi_pll_reconfig_cdc_m0_write                             (phi_pll_reconfig_cdc_m0_write),                                    //                                                    .write
		.phi_pll_reconfig_cdc_m0_writedata                         (phi_pll_reconfig_cdc_m0_writedata),                                //                                                    .writedata
		.phi_pll_reconfig_cdc_m0_debugaccess                       (phi_pll_reconfig_cdc_m0_debugaccess),                              //                                                    .debugaccess
		.phi_pll_reconfig_mgmt_avalon_slave_address                (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_address),     //                  phi_pll_reconfig_mgmt_avalon_slave.address
		.phi_pll_reconfig_mgmt_avalon_slave_write                  (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_write),       //                                                    .write
		.phi_pll_reconfig_mgmt_avalon_slave_read                   (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_read),        //                                                    .read
		.phi_pll_reconfig_mgmt_avalon_slave_readdata               (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_readdata),    //                                                    .readdata
		.phi_pll_reconfig_mgmt_avalon_slave_writedata              (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_writedata),   //                                                    .writedata
		.phi_pll_reconfig_mgmt_avalon_slave_waitrequest            (mm_interconnect_7_phi_pll_reconfig_mgmt_avalon_slave_waitrequest)  //                                                    .waitrequest
	);

	soc_system_mm_interconnect_8 mm_interconnect_8 (
		.shell_pll_outclk0_clk                                              (shell_pll_outclk0_clk),                               //                                            shell_pll_outclk0.clk
		.DMA_to_SDRAM_reset_n_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                      //                   DMA_to_SDRAM_reset_n_reset_bridge_in_reset.reset
		.hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_010_reset_out_reset),                  // hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.DMA_to_SDRAM_mm_write_address                                      (dma_to_sdram_mm_write_address),                       //                                        DMA_to_SDRAM_mm_write.address
		.DMA_to_SDRAM_mm_write_waitrequest                                  (dma_to_sdram_mm_write_waitrequest),                   //                                                             .waitrequest
		.DMA_to_SDRAM_mm_write_burstcount                                   (dma_to_sdram_mm_write_burstcount),                    //                                                             .burstcount
		.DMA_to_SDRAM_mm_write_byteenable                                   (dma_to_sdram_mm_write_byteenable),                    //                                                             .byteenable
		.DMA_to_SDRAM_mm_write_write                                        (dma_to_sdram_mm_write_write),                         //                                                             .write
		.DMA_to_SDRAM_mm_write_writedata                                    (dma_to_sdram_mm_write_writedata),                     //                                                             .writedata
		.hps_0_f2h_sdram0_data_address                                      (mm_interconnect_8_hps_0_f2h_sdram0_data_address),     //                                        hps_0_f2h_sdram0_data.address
		.hps_0_f2h_sdram0_data_write                                        (mm_interconnect_8_hps_0_f2h_sdram0_data_write),       //                                                             .write
		.hps_0_f2h_sdram0_data_writedata                                    (mm_interconnect_8_hps_0_f2h_sdram0_data_writedata),   //                                                             .writedata
		.hps_0_f2h_sdram0_data_burstcount                                   (mm_interconnect_8_hps_0_f2h_sdram0_data_burstcount),  //                                                             .burstcount
		.hps_0_f2h_sdram0_data_byteenable                                   (mm_interconnect_8_hps_0_f2h_sdram0_data_byteenable),  //                                                             .byteenable
		.hps_0_f2h_sdram0_data_waitrequest                                  (mm_interconnect_8_hps_0_f2h_sdram0_data_waitrequest)  //                                                             .waitrequest
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),         // reset_in1.reset
		.clk            (shell_pll_outclk0_clk),          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),               // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),               // reset_in1.reset
		.reset_in2      (aes_reset_controller_reset_out_reset), // reset_in2.reset
		.clk            (shell_pll_outclk1_clk),                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),             // reset_in1.reset
		.clk            (shell_pll_outclk1_clk),              //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),             // reset_in1.reset
		.clk            (theta_clks_outclk0_clk),             //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~hps_0_h2f_reset_reset),               // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),               // reset_in1.reset
		.reset_in2      (phi_pll_reset_bridge_reset_out_reset), // reset_in2.reset
		.clk            (),                                     //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),             // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~hps_0_h2f_reset_reset),              // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),              // reset_in1.reset
		.reset_in2      (reset_bridge_launch_reset_out_reset), // reset_in2.reset
		.clk            (theta_clks_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),             // reset_in1.reset
		.reset_in2      (reset_bridge_shell_reset_out_reset), // reset_in2.reset
		.clk            (shell_pll_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),             // reset_in1.reset
		.reset_in2      (reset_bridge_capt_reset_out_reset),  // reset_in2.reset
		.clk            (theta_clks_outclk1_clk),             //       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_009 (
		.reset_in0      (~hps_0_h2f_reset_reset),                 // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),                 // reset_in1.reset
		.reset_in2      (theta_pll_reset_bridge_reset_out_reset), // reset_in2.reset
		.clk            (),                                       //       clk.clk
		.reset_out      (rst_controller_009_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_010 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (shell_pll_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_010_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
